`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FZnznUM6enUuX8LHrmo+1QyUeb96vezNQRp68KOCqOMQ9iwbSXXOvetLb3EC9S643dn60YqNxe8/
0c2OvYsjeQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
hfc3XU4xygrUFpaR8EfxTI+/j7BnAOzrnZcvBSwlkwPQYvBrQfGgpdwiBlnz20Zchc+aAkzLpAIF
QmjRsMorikmvOaYqDn5WQOy1VgqlLGadLNMYRnFH5nT9Gcpz0FzkeAT78YFFrGS6G/DUVp+r5PcB
OMjUdqQidxkK/oQ4Thg=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
tVL2z7by75Gq/y3sUJL4Hc+ngOqWLVmGJp/XY96qWoQUlT3y8ARNPHsxkg/gaZihxJ/pt8H0JiSP
k2D/Gx08fh5DHh+S99yuJtFf/0o8b2GUVbvtm9dGd3w+BxOsSaGrZcvrhvggtp6hiY1VsCjFT/uC
bcDmuDzp6TDmT7whbT0zxHLreK7cG95EjFO95ZtxEXW8jDLdIM9XnOk7UO3kUj9A/QbFaQXaidAS
Mz0oL0mGFHIYX0+exSoZY0gJ/naPxg3krgBPglnK31oY7aiP34aBNud7LpgSh3M2VZa4vf+MPR6N
iNqklwoz2Kq0StpXqxp03adA6wbXKyVCmv6iDA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qTU67hrGyd+x5voTPsYZXqJs+aUWKRT9UWUWQeCQVcYrGTFQhXpebEPnBwaCDwKIS06zXDsyh6JY
pTKz5LCv166G+B9YJnYVeMOAOfI71Ftxav7Gy4FFLmYrCb+u79HXQQaGtPMqosjvtVxuXpQJEejp
//X0QpkNuL47gnNEOUuS9D148aWnjLZioSHm9IWaVdPL2cJ7F6XEaVRupnB0nFdJReEAA0glnSld
r5VmJ+ousm/1QA8DaOYR4nMFhY98kKqzXrrXEdxmfqa8xtpHMxmd7W3fcuc8AqL5/GXoeRctLF+/
wlBjzvJHvF01XXNJj1TfNHa10ApLYTCJjDmlDA==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lkiXMKuo1I88UDCCmVVp/P4UQ0BWT9NaPiMJRFJAR9Xic78U/346s2tIqCVlu6kJO8/ypic4dFx1
OH9j9sW41RoUj6rwEl8cE78E8gf6UChbTB3UtNGZonM0lb3vEy1B1aWfS8n1va8WUb+k7/MjhhaE
R1/r6A2+WEAO50rJkxikmAgoV0vJdVWwwJxOWqk7QW+aFBks9VJdfNwr8+ct1fmW5USwa+sOl+z6
WC7vOIUoWVQrSfCzYtLJJu9pM4xgaa+dkJsAclkOsqCe5AWNgxKQZ8ix2wr85CFj3Mmb0ZEM+vBo
ViuHNXCW6dY1u3oiWoTvshu0AemSX4eGpOl1eA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fTfxFy50qATOYlLe9Ka9qyCpD1L+4pOu+reEsUNerk5p3eTV404ecPoEv1b2OqL6cNEfKTpoGZB0
glwHpa9CWM/TvirnG9bO2Ll0dzpT2EDFZTTcf4NhfHOxQgb4fBGG7uXIoR31FjJspEl0s4uOYATP
FLG8PBcWON6hGwTjMXs=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
V0qwZink2QcbN5wPywJMYkiwdFu1zDg4oT1fokHYVonExoBJycsM92paTunsZndIg4KzuB7WjrN3
4TdLM1Kr4I62nnI21zKDbKN9mh3GI5nkPXi792eneAddudiaffWtmvmD3zeaR6ESYU5TU/H8Zgg1
1cbIpz/SAeBEjPeWAPRMxvQDrCKOQJI4dADl4+qkJ8nww7H1Jb75IjxtEDCbR7nxFvd3ElTz2YdT
aSWHFJ7oQeYQNero6pDreMT7AcZq46DacgOSgOPHxpcriNBQlNIMP9RiEGiuFCOVXnWIDHMA0p6O
xJdntDYu0lzDcQdaYcSXl7ZzIK5JANHagtb2uA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 70416)
`pragma protect data_block
sBaUPNaCeY8MrRsb8lX8n0uWrlftHIGAi841LNoaj7t9Y+7eThuU7qrQqrOyP0B+n3KQi9hZM/Ob
HlMvqOaUhzrQiWjw+6q85JiiTNDN8P8Ma4bvA4ml6R+UxyvuV3QAyTgKBg3a4sts9bZLHIKKOlHA
lYvjbUOEjr6PaIAsSO66LhS5UhtGOfGS1v5ESkKaXEZk27ZjqLOmSn6mtKxF9TRcuun5+cY4UaHA
vKoejBXQyFNsbOHoRrJNdUk62gmeK/1oVjS5gYqFqJ6m35i86q2QQwbBoOR9TX66WG6BEyYBM2Yl
Il0TxG+Tj/PsxmGb5M41kLiAQNCmZyocc6Vr6wVvK+sEwcfUdh1u8eKtSmvnU/uYq8Cnbm4Da7ur
xa/bJGOqF1sj1zkIi9fKMLA5mNV1bKMNKya/2/gsGaXUJ27CAcj4+Yy1F1Q9PpS9IWrGYdFg8k7s
vbIHP2Nakh/N2V5oqY6XWSaBRNfKKjQZOuaeOxN0lL/FSQ518BNmboFiXNmjB6PPur9LZG8y20Tb
OLkKoGubCmwLlJgQzYL+Qs51Zyp4waRt1IMMC5EAHW7SV8uHxlWLubW1UUwZjzgfjQKmXPQnkT9k
Wh/WyU5BcKPxL6hQMuN1hN43jB6Yjr1vNFNbyeKpT3eBNoTBPeVE0u5IEi/rPwES2LBILCEGxEL7
gnNZ6usU/K2UbtrA/5rZsDQ1EeV1IP0zDr0J+9wGjdamxinS3FfwWur7aePwmTaxTlmFgt3uhowe
P5adaHY/o7ZPlRH64mbHsri333LfSuaD7moBm5oOOZ8Up0DJzYTA5/CWfthe9H5DhWZnTFwMoxQB
0c6WTeZrzDH2E98TQIxN7W7b9cjaPUDAoHhxhjIu0PA5JzGTIXuWLcz2pQygfs7BZiRiUgxhlqu2
ULPCTiuirz3JymmBVnyTQVNFwBqwm3PTQReKJ90RAiwgoo0v8XEMj7ec7usjIKkEk7d8cwXFuVlm
7lHQqmwnRyZdqcmfl+EiUq3uXgD/mCryU6TbfqFBp/gUKcn9+dC5aOs+D04mDmy4UlWsiqGLFsKJ
kNEhpAQDnUtToF+OtVISOohWp3dRpabTJjT7bzcBa7xu0xwaDCf+LtXWc+imhYnPwtTcS874YQJB
AScqqnNbun9AJoL5JyjdimKdv96qIIORWMiTN6mS6rXZVVxFIvKaaY6iuo/1q0p52Vnrl2w5hd8z
A+Ye3lLrMIhstaTjsHYfcKnFcIoWVGNRaVAgVYnXzhG4HMWF5ZX5M8hXaHFUxDvtewFLmG+jPLJo
U83mW+Eeb0lDS4tq+4gZ1eB5DQAekQYWpvPWRG9IWi7m4PJjgenoP4c+U9hlhkasbosyXyH7H4RA
4rbGnXwyvqz3UUcD0hhFQ9w/lRphx93/KbY+HeGPNjZn/cZMh7c+qC/tzWspHZWHdK/fAhWFW4h4
Js/iNdprtqtf+7+qxA+Z5X4qB1CdMs9abNiic8kul0izXZOWI6CFiV2TzUaJGLCQOwf9BOjSt+nd
YkwoMw6yuXwhDqg/Pd+ouqZmXW9bqfnqCBBNIiy6lL2rF2DwneNpqUtVElVJVdcjSzYEzrstmQXK
euXOPBPaKYcYuSdUOEUyN+JeRRHSgjxW/1ZXbg+5tAE8dinvYZL0EQkaOBF1ql8V4RsmOUpck9hH
gu/oJZYtogMG3KBVHxFrZ6T9vj8OaVHga7JfCsYOOpqf7TiYqpKnUvhj2Fq5Br5bU9ZtRH8d8rmN
jnXPPEupQr6DM8r7koqaBnEzLShNsfbzpyqgPdq0SvV3IdyJFpYSQAn6lq1n8bjv3nS3g/WRWZUI
0CHkGgCvWD3hlqPOxD6f5bKi8NEThpQfaPZToZQN96K7kaX+wFe3EWkpiNUnMEP/Hal159ODJdNL
jqMaaqMVxxx5vPb+8yP5i3bYQWGkO3FYHJy8o7BQ/MFwQ+H5ioSAM2rcI/Fud99S5Dzm0o2//a21
IeIjI+FZSfNL0GCDgv4boCYWceVFiVLb0/CDUAVnmDR2P9t+L+X2pwo3XmRB19HxaexgiErynRWg
y+jsjs1w8qdP1OxbThAr5BLRi79hNILSeL2RErpiPmdYEWEglEUmQrLU0qSJ8JXwziT/4A6Taa2o
eBSSN/UOHgUANYs7fFkVSSO9aMQ6lS6HFIbxLyPbkL9vOuSLwaWmgL6yy1bW0BNqe5Aq1fb0D6sN
ZUJeug8XTf+bLXeZIqySjsJyHP4HBqSV5zR/j5AmnAQ+/38F3EYajut/HQzio1uxwcJeZa1B8Ib7
TMcMQC65mPaD6oybi49EfaQxICkpb7oIllLdBkZLib5FYdB7B0FHOQ7zKwH6hM6Oc00u+1djaywb
D8nSmS/rNsfo5knvFaHQHcT+0Chk/bzElkbcduyYqBEat/8wE7aVVipu6L8DhIt4T0BQJH6Eh5Hd
yVbnbk3kxMkM3o/ENSCt5ThkNm/J5EGJVga5frgG9zpinATD10ccX1WghnhV+6FuydiVq8bQ0//l
IaRs+QebY/Y2Nt5VZVMRGzsLMUwGTqHYDvEd61sUEkz4aICDEncICoyeNUAVMEdRMY0sJ0Z9VhXa
+dSDLA4Smnr4akb3835GbqyZyRqICgKWc9aRc2bZoEraUjJO6qMJV5aZbzK+00yx4nW5XinA0uvc
TEYZIDFdDQhv3bgRXoPf9hHzJcntPd65bHgcqfpK8FeIoegGuX763hem3NUURwtGc8G4bsQl56im
/YuX6tMbUjbKscZVZ2riVskjRg/9B/kbuXdigOB37AbWAFCt27VEuhL3HI/E4g15cuvlD29TaV9r
7QswmPZLajGGDUVY2vLBENVflz3oq7gIup6BxQbb7MxtkAmmCg8y1WKBCiSrWguD47dyJP4QvTzQ
5493xqU8djUP/fnvg+Lcp2kQmpbTs4P8stBTIplaDDa/SAzhSK/yAIBKnAOvm4SBhRUfTdlaRLDB
ptzXwcxwsECP3cjExJWX0hj+p/+vGXoLZppP0ZFxGbA+FSanRM0MgVwcoA7/+G710J6MgnMhmvAe
MsLZ0DUC0mER6vbH1O9y/AOhFOfIwo7vDIE6i+coSB7SBhZp3TGkmF3Y0J20wuOFrrj0xVtGgdSZ
hOkVL4fN86XOMRMdKHUJrq5h/h8MV0hrvh5fXbYu1B3A7X+sSiKQ4HUw/aM3xkhmBHm15VVO3Cv4
MEhQyqWvy0cawpyaU+hsTTO/S9Jn5+XSmrkY4OyuTUOKEmYgs5xMwG5N/Zx5M3W3wuOv9SjtdPZi
u+gatP9lTKgs+j6CgVXX29tqaHdu3M2ZlnhyPI/TqPzQMvhlL34cXhJPTUmDnFFK4IzxPfU/ylQg
grqCi5ksu2kLCmaqq5w321SPozKL3O/516irFjqVKpC+/SnjUQvsnLNnIye9B4pF/UyRd9sZp4rd
PaG7HT9djAwll0GhLWg+QJj5xk/YlBirEOxaxZRx/4cMrZ2UTaQjunAhoE2pekyA/kPtz+zGow1A
WElVAzF0ogtNLWYeEi7/RtLKhe8e0c5LdaSS543GiGh9k2uTNo9v3d0TvbDhW1bNuBJqEFY2MUaN
rlDUhbRXgZHDk/aS0BpyrFwVGHYokiOXtJFH8yhmEfoMesHEk3lv+Sq1WDhwkkD9ya6JFMXGVMiG
GO9+zjYrIVUyIv1kQdnVCQ/vxssREgt77DSGF7wPYT3rRlkg6X2xmh+CEGOUfvCw5XHMKKpzT7NM
TFC2k/SCoFWyEuLmRfq0nY3L+G95Ats5kuZ59UCDCvaiO0hdOe64seKBYlVdlv6hwhwv/jI0UTwk
Ae3S7btQW8FmVgAFMkaf97Kgk9q6gTxMIlXFDAzWnhz6m48aprkBz4gb/wHFzxP7XzQ+Va8LdF90
P0CkxHiXWwyouk9dLKNQgzBxoh/f2j7DuyRLFljdZ8i785Dh9Zwoa/O2yBBKCrpe66Nz+uCRVo9o
xriRHJPp5H2Xc0kdSX3hj5d4ulU++8jsTZ/Q3tHA55WMZwPRzHSrTJO3oadIxD1piI9gLw73zcZF
DojyDVQ1O8gDTwsCpzjcQMLfu3qi5ECK7sdj6BJIoMCiTiI1n4QtbGLjUrGWogZJpASXM9dS5iBf
NSSVOeuAa4ssRV8cuZwGec+4zGoTuQkAwkD1EmklHOrZbnLG3ELeAZeFEFjAiSUwC8ZrXs2BBMmO
KWesBdlTGIDpzrEXCgl+g4q2mI5xOURvbNPb1Eu1Ew35WU85WknvsGVIb+NLC9w/18Xlvo1J7oyC
1nJ948h36CTPvdBVQ/aAKcmjQaBxBxB9ubvmSTN5GxT4Q/Ptx366/M5UY47rd0RgMkUjpZ5QMMH6
+Sjv7Yhi5o3jrHMzy2CS1TfDYABt0BVFrl9rNWAjSYBRFVMG15L+ak13S/lbp5tfbG21Ow6OZM8j
//YaH8nK0LDo3wdF9ciuUnPsRf9nQnsZVUFcRQb7vuTGz3pIUEUJt1HL5MTWQ6CKFgCOsJZ7A9oO
wa1KQKAbDGoKW3v46tgYGJiXeuN7prP5clx0zmUAKTmcINl1RJ4OobH3tR1jgl7+Wv9y/TuggKIr
0s7KB+Ryo70AujiKHuOoKTLBsrQk1a4pcaJa9975s2nb56tMxA3yXaMcwK5SUgMMJj6P5DA1hv9j
E8X/8xYogltxPMkec3DmHed4xQH9tdyOIN7PuNzuuwnPvRcGV/UjBKZrtgixpfSJAgzfgIRaiKwM
2KHBvbJ4aCnZaFl0gaiZzSl8GJTUIWIlbVFrTbpgYd/lmrvrmckR/Gk4F6D/ibbOqHlZkkhcoZHu
Nj/1uOWw4ZMyhmwPAKCFo2Su3ymPl8QjYV5V0+/Q1bKwGyBg6I/YM3/zraEE1TwQFyjvzpsCAtnf
aTPgFxl2y1ShUw4H3mGcbk4UyxJgschl0W86lh0zV0mgzdCG05pFfHyOhd+2yc7/kHT4FzDEy1Um
rc3UapdQZLtvV5V/If2QtjvZvpG84H7Py18R53eGogqb07dDRdvUNVvYOMi1zEhqyRzYwoGXAjQy
r4jWZ+pciI75xYCEriANq0jVZuKsdxB1vtvDV2gsxq9qQ1kdbDPh6AnMQFxuu1xxQcLDNQdCKIWD
CLF9c4YWTVBpm69bJYOoOgfSlcEiAKHd7M64F0lWr+7yaCskm35JkctJT0LfxbhWh3HM4oiaAhtp
2PZlKo1qFEL0HoJu9R7kSBoeVFkxCvRqD1LCJZWpuOqh4APyookY6MjQFYr4Fce+wl5mQKbpLbSE
C9AqsIa1VWloL4nBK28PgqhZAqNRn5vSoCIMIiMFjNigCFn9T/LG6xxV0Dk32P5DTYGBYSYguUoS
CjWq0NuH+a9D8tllOF3+9AciowrNT2F23NheCjCEU6GH6cjaDFVu4qtL8Mzj3+35mZH+qtwM6Hqf
VYo+dEZkNHTrkBcKthQZWtTXiFCyDO7nEpeKoGY45/ipvADCPpvnm9ezRss7wocaigyV6hbA20sk
wF0GPaubMJCs14tABYa/vUkupnsWSu2H5hnZ3XXgk9qdYrMx0a4JBGwtECiWsfZ1Gsxx4DmILW8v
Z2LoLDezpYsHAO5x839W0kEer1FaPoA057KM8WZ5VpcvXfLUsqZCtuU6GPoNLGGYid2nFAUfFK9v
c6k0q2OR/5zKw4/lLb+DEm40q8nOruMruoi296qJakzai3/drmqIGZMtMCEWgC+DoRPG3MVnMbg8
mO7Df9dZzip+Q7P/95j6fVy79lya5EgQRL3f6pXZpqwnXbqJcrvMZcI/BwLTXaNpGmIJkmJr9jqC
yiYNo7ziGiarfmLHG1+uG1MPI2IiC1RS1T+Tk2yyYKx1RhAaHjy1lwBWrcTVTxcKE/IunMPfPBBs
QWeLvnmN9kZE32Ey63QU5HSZuye4/VttHaO0vzh40V3L7gwcALlwXZJUYJ6DYHuSST2GKbBs7CRU
AmesTkfyJL+B8husXyC7KdVkHUM43Er5RD2mc66ZoWGDi/4QyYlsnayz0uCrcGqtvfeV51ElmS14
5LrkSLy7VlmyxIbw7p3qzBiJmzQ36tvelub+JK3mWd0DQXTx7/uvvYmMU1vcJxGmuWJ3D7L0Wubm
QD4NpsRMTfJNVLEC7lACCztWfBjk+Mkuf7SM6CSv+21OV3tMlo9W2AkFLGEW15b3AgaF62SfPrc7
Rh2vsdgKfrK+fhMMGmMnjeQIIVRJNQtuO4HDq4G3uu9+SxVB+i/gel17I4yaYdJtBHj8gLXvhtUo
LIaZTrOQGhZNb6yKltVdiW1xUR/Mnd0b/pVXvMcaWvq0Y7OXyLfhK1GleyFCWnTI7OlTruiSXRSE
KlhqmPR0lYlV4s1TqbSpbMsHINZbON4UnR801CNb5Ul85C7XnyixZvaXss6aYridnMg+1Eu5CvxI
8FwKU9ysj+ySYEKLI2K5xE+a99vCCRUNKRd7PUQUDnqzy+S1A4ok+6zO4G10O1PqmTq2E6NuCm9m
2yJSZ7pye8t/PryCL94Ewuaa8sVS2aIHPP9j42NDwPHtDhNU3BoqmHNVR81DNI4SeYy49tBce1qy
VU/CYO1gzcA+Tfc8Fp46Xa0KpO5+bntLb5FiAQKmR+5GZX0gh5O8Id2rfkORfmstzzQj7ghY5MME
a8ZpT53wMvoHqpf99oChLO606gIdW1XY7cZ7eOJL9p0+kUHJf34VMS2GPzRz9R8ick1zfv4frmul
LBzx/5Gq8P4GThpVfousk1nrc+ZEDPVevzEJyMqsJEOMVN5DiNzOHxLpvD1VYP2E2iqjps5Ri7vz
6PKdskIRo+cajZroj3uhaFV5nl/cBVX3Zj6HDMBA2rQDEg3cxSMHNIRyhiSB0OnNcyk2Kdxhjo5Z
RoYDfBpV/y6GmP4k0AAKoXpbhGWWr9QKHc8FLRuzpbGIBZYo6iF7nx+JRC3a7EeRa0ABVTnGBHld
dkFlZzCVUbITPgIdLt4386CxZhclUjYzTbdy3jsxRYOeG95BlIrQ8CmV0zUBtv43rJepFRQJoxog
p1ocdf574OSfH+yj8KZEMqBjtvia6XSoICcr9g2mZ7AcKtE2JxT/z1wLm7BUaJISU03qdqaJBez0
DDMU0iMWR/wPsn9y8j4mkdMGmUBMi1m1yaa3e91Cl+SuB083ud2wtdQjCGKCj45R792C3ukdEoQL
fZjP5kIpPfvO0p9RtlJqyLULIE2n+Fu9VLl2OPaV1xg08ce4HuhlzW8BlPQo+OkEgb3RwzF6prRa
bmUxk6rHNsab/aqXchvgFXMQFleT9PhDyAdUyNaB2Rm3SPATzRbU0443cZGU9RRLv+etYN7/AVF7
CPbb2l/oY0o+tpDBU9p9PRem1hCfQVK4tlrn159RZSyiAaxpCPKxIg69N3ASxr1f5mNKwmmSLQhW
ngf8eHDOy15y5uAT8sqv/iPLfxw7FMYmGZZm2zKKfV59hYiH882R1UuwCQ5+7DGQdk91WGOYf7G5
w58DjEGcGHgYpxtS1eack1Wm4ByuDNsIk5iV140RqYtHWbaZXDuYHbdQGqXqQ5XohVa5Xh4We5N9
IXUA+X7KC5CHE5w/BWzQtzcg+IE+53qY/2VQTD6m89SVBATs3nZL8sxTu8mJalrllJrmnV8Hrd2t
kZyMkqLxa3fug7Dit8akPJVCI0gjbOfQ8G5R1T/SphdT784U6iviW7DFKdINM76QPdjW7LHNxrDi
o1gZPT5RnW5USbue0YIpbZk1ALPQAbtKWCoUqJfSnJobJ9jVAfmZfIXCxk1UIwO0NJ+PeIsAoxtg
djq2MPVQ79LdTsvs/X7NjYOzTCzuBQuCt54PfYrKQqgBLF8eqycSMLgxz+RMDHR0yKxfdmy3laG8
+Kib/q5YS7is5kqQjisXFjlhoDfAJyhhswPw/FVYWJ7tQUD0TIgumiQUzjaBlS79oJuxGQersNhh
fMKp6LDSv/uYbNFUHKVArRuZi8VXaljlOlOaKlXXYT2ND8VFzs5Ac5dHRCvDewtpzmIqfcixcF1Y
LMVfbU3AmibtFJmCQwlc59Bw1S4nKyjcJZda6GZQRs5wK1yRGBwuzidVrVJeGKsmO4XpbyYZCWo9
u4LtxsQMxZVuzsgfu0vOhnGNQpAxDF1INutUfYpLAZTKTCtH6X5nKY/N+0QJ3GU0gixMkORIMXX9
W+0cJBywfuY/Kwf6DrdCe9HiOFJXHvWNu9hMFvqNMF6uoD+/IUTjDFRxLsCVETbqcywJso0EHNwW
klJoBvjO0fRHElGiFfATC6/X6A5PwznP8n908/700oiMtwoVbf0gsqtUknkbNk5axabm9m/rkoV7
a0e2bBTdv93x2h9zUAICJNagZPNZU4VyNIIOHOLtzgwN8yVcTdYI+o0qDwEGetKbUFpdYUkSkS9o
zwURWxBnvQMgYwZKkcHeK5fNfMEVFlIPCKYtOx1e7GBiU1iEXO9Q5+iyKt97ne2rAxneOlDNDhL4
YyxVur3ivq7EYxKgXdGVwBQ10AaZJFLUFKSOZ8iYas9ApTKib7yn0zwzzqadSuOknV/1S2F2Nqan
GWcV9hMCAvZWla58QHpi6A7w+qPncLRcfFqj5NU/lTbjJnuM/0mejdk94Yehd7Q1uQd64FkdXzMf
mQynMnEmLKZEtS24ntrLp6dTsGnhScUPyXY8hc1DKpjEGeQaFaaxeUANlf8ToYOtsHQmjZoaI8rY
24sHuh4bsjSnPW+YATgNvM7L17wWlLpPcNKcO1y+wCyTqes7imNFmtruC+UqHgBtnOSsPYi+4IGu
2+/T5gQt9VUIMKmiHB04Lmh8w4vziAHYTEKhWiE5OXNsNty0GKsxXayzy0w9UTItEC+klXbwkRHd
rsjzIvPnxvUIHjL15ZWAlP/Vh0MAcHmq375wi+MhldX34ic/jN6PUVy7kXpxMoolqnC0C6NGdHUC
SXc37gQ22Ah5Jr9HPUsmFC0hZScmdJUPHbmO3jPv+lizv9DJ+mik22rpmNa7vtGOwIsWPYvWPcnN
h0rb1Z8NzGoFdm3dvJMlqi4OEytxqBegOd5v/WjUdiIYZLNwAmhJOCO5OjTs+j+nNfvj0lb9pzGq
k/agT92FGxiKlH6wS94TZ5Ihamg1Zx7lLQfidl4h82m+RzucZXSNViw3SkmDHmbvRZZzeP1AdP71
gUunpoayt/BiVytXMZhJ6kd67JlYLPuUpccUq9llF9/2Y8ad7h8zdW3eretlbt4hy6Bu8LldprZb
TELX4yy/IRONK5s5sgflcngxX64EM2eAWxxYQRQ8GtRA3hjo5ZcgBIXNzvkmRW/Z8TJWXCV2lSwB
BksHMBKHyqALvBMxJJ9FeHkfgo+gD9fWBG/DJXO3WgBbTBsl2suAPMapaunYQ9kKuDWK1p2v8Kjh
/iAi9Lv+BXiZDWsUvztZIkmOa1tUZZ/fOweJSWTyKebAf8Xs4KiGn26INaFR+ZiIRF6DKcv3sni9
+XWNN3hE0YZ+eHXjKfbP1RP1fMbDfYALgT+CpyJlYxyG5NGXMfuRozDM9Uc94P/hHS5RwETuZKzo
rW2t6wBkUjpkSIURw4UjEq8EI1pdWUVV9iko6NB4yTPOJk0ii02ik8SUVyc8B4RUNsnv0r5AxZF6
0YICyPbxhs0NbtiOvQSvcXWdKpLKBsdERo9jNr2d18o2D/coSVOoL8ke+vhH02vD2Jd0vrZs+z27
RnY9zKapMNgSOrlnlY4x3iEd3hVBTd3JCc0wrwB3Y0eQlwPO9L/CB5+K4ZNZgf1OGN75XmbICoLN
w9IIfWoTif/fzBK1CF06lhu8sXWS1IhJO/IoNJPfk3rFeKR4lp3qvPx7qdq3JydA8ufCTcZuuKb+
SXtBme6VLM3haQPI+mj1Ye/0JWds4rPVmhj82KkQuZXDG1QlqX+ObayUiQ1OwMK7L81ViVLFJKxo
9HyfX8MW/XyoIVA7cWtqrn+U2DHtk7sy0ejbc+UI1c5+0ryjepFE6m17IYcFt33mr7unwH27SV5A
fw7Oq0EnGu8R0RlihVMLyspcgHxzvwbUqBTy01xjZlUymrJ9WgVDl2Ek3BCGHUhAq2IwKJvZ5GPk
APibZQnxKd536VJ+znvoSUiaDIvnOFW+EOiFMsYF5+9WqW6evhcv4LMUpuPrI/tC0OVYEnPbjB9G
HEma7Dx8exATmtXOspZdR5G4FYHKKD3ENOaUMjU7fW4Ndi8k1Iyj6yzsCSkSBpT3R6Cs6GX2ZAgy
zL1/CLgU+6DrSHoesfzkVJDWUZtDR8h8CGj9hkATqg9aYpSMiwo4CO0zIvY0bfIQWKgO+Tw+E0A3
NBl7WQnvtgl48862hPFI344hpg3QU7qoMs8c4RYWXfY6VKmq56Y5Vpm0HiPZ7qbi7Emsz2pDcf9H
yzP7s6p7G/Grk6m3981R79FxBSeg5KxxBEiwhPpvX1zSgXNBunKBv/S8UPVxoKFGIkumXyTcpL0G
xU6BJAGR5HtG0hF70jRoVkEt65Ns8KTVl4mhsXhngZAERZjcZI7eHbeV0jy9TRAwzNZb7RZKwn7a
oUtGMTlfHqO1Ej/2dh3ngbKZTIx/3zuyenenLDmiRN/mLqNyXrhqs0Xgxs0xM0tQ+hioNV628yOj
XmJhaJxZacO5SwbE30l/GqALgK95toHOjm+QHHMv1qHwf5tktWI3WPEMv9umB6uBNqKEQgRvGskY
tu0rkB2hjashkPXA22emzXvkQbwgbRNl1/I3fbersEOvj+Ujw/fGXsYZSlOhR0/pWz0a86fDUhYF
TOfxtriR3q2HT5Pr7vzOR/fcuaMAAc+av1k4PARBf17Bulf7rfxlBum2pd9ZFqFKJWIJPjmJeNuQ
eFKfjfVPY1glDRMbvCtBdOJwTzNHZdDJMVrODETyJdJ6n8lYzBBn1dDJbf0Rov4tr+8lQzs7GFJa
y+Oh56Snf5yI2SZTBP2fISQd7E/705nc6tqgitLiCaI0ByMJmbjucVLeUSAhwosjDhO1XS3/5VxA
XqbmaDsthVjSMuhAv7fA2HFeiDZ/Fp2CwJjoFvsMsdukkWDmEqIa4IuWaoU12P6CpzDrqbYFt1li
HBM+YaYNIWmxb6nOomjF9T7hkwJkQszBiPc7fxMISb8iOwr7cUlqIDSVRpYzd6D0sYUfrDNz1Qbf
p67T1+cUk4oLdI//lRt1cNl2et9G7lME6+sehSdvJs+mg+WrfmIXq148UNH+kIewdBa0wkwTqG9r
GmEBn+B+iKnjvN9te1Zu9J8JBjKjga/kCwEKbiJHHX/lUhmMve40m35/707QHpK1Hk16I+nwUWQz
P0ad6C36wyM0k178yoDSaXSi7jOTopnI4gH9PLbZQKzs82dOdlw70VtwJXlVfQzUtBTduKpeqzKF
Mm8ALepAH3NbfkITzoPCSQy91BmzvIfT/lsgUVXsmT3x1UUkdb0ZSMIrnjt1U09bs3kmYyfzTc56
RiiBsdbPr4l0jF7tZom+Q2rfoOeEioOWRU8y4FkahiONXE6srthVh1Te2r6HcX1MtO6r3dvFr3tn
Q4Bn0XEQ1J7h5i2jga7atT8klYAXHD7XqcDRyIWXsc3xU/X204rlGxLFFwGwnmIB05jVR2suIzJK
m6s4SRgmjq+4Mpr3mL6y5EK9gOal2wG6gsPMv9KfWTKpcndA2JI+/wxVGeXTI9aG4w9tM7upFDTA
SLdOi6EERk81tPFuklZK64dGxiaV/ADAAa5+sBPKkcQhbh8wjHmeLfS3sVd1u94UH8Qle1LpkGKP
BVLVnC8MMdCodUDY5bqGTcAdgbDBeaUqJOx6GiHAhAy2tjE25ywXLydUN/kjO6MpyH3L5n1NHoEx
6HzygCxFNUrSgOs6rzmOCclbyWyiUYTv5M0E6zC4pChLVc8vK2MdApqHSVFoGXtZBR4mkQ5BN9o2
cVDSjVCeNHkRNymbF/uQQihey+qzmRHhVLkcd9I8EvKZoYFgVJ0o5adyIim6sZ7wVAzyBd64eADw
v7mAECpIJi4iYjvnRI04RMfcUFpeEcLnUbrqLqboqNvqOTCxt2ZW9vdfax8+XdVvaWBGPexP9P9o
mL6QvLnUXkZYGqgMSFL/pSOGyEIrZqHKFCno9idXdvNvCGM2c0gF8q7INmMcYU4ZqbEAJs25rApB
vPFR8yDhFfR8cJwjleojkK03rbPVTyNhDGSNNWw48drSrh98Jg403WpTfBE1JIjVUcsh+3AUO0SI
svPlibEpTmn5T0bQJ5BPUItm8eE1ynJlU9ijBes+OQBXwscis78TD6HPO0mYs2a0VG3WjX2XRxxg
qep1krd3XQBsEFXf7NL/fINhTTG3bpurkXHhuENgAyYTchcvP/YSOovx3sLc7SfjbhKiz9euA+F2
CFGCDBhmnNec1c1I7MAYppfc1PmMbOCsKTP7AffwOv9e1yPgBHkiUuY6ohcJrumYvFyX/zO3q4gT
auf2tRm+qHE+xxdc3pJ2Z07/bVyKokGNO1VAv8lXd4amD/V+6XrPsGM5K8qqkkNodORSLT0aC+fd
pennWE47n03+Vt9CNvcc2I91Aoz38gLKhPQqnJ1OSKqfDJrQEPRSngMt6PRRVmdFO/zY2yabbvnt
SX8on8PPhIPEgUs6upjxmhU7dYPjtIO7taIDEEfqWHcP0tgC/FTYeLqsb2kAIJYOhGxgQm2yuHbS
FYXLuRtpoeO54DPYHhLcAdgJxA0qt1prCNW8/vJA81lULqmJSLHiWjTjUBlvpsNzydp4xutd3jxK
VUyNqPLNyeTIppPiKLaD58niKiYRB7SNHVwitcK8Logk+THOyFgJVdJ/3VVwNvi5fhdAbRx0AejD
a1AFEh559THnYDoWAbWIji7SJ8IE584aRf5roqNwD2ot43dxybXWQ5rxmO9bQvnxfd4WF67a6DNK
/NRICdkOUvq03/sX97PXgpc0wNGHA3kq8toe2lPsC3PfjnreDLHHp+bFDYq9+x1lbmPEGR9fQxKX
pn4n3/lSoD6jhrIj4/ruKdLCw/MnzrCSYcVG/2Em1255QDTtQzJT1bvoXh6xE2eqccXZOgGKj9+b
lSfT+CVnr9yd9VaE8Hay4Gn6jQ1zazQv4QIG3aTrUBcdGW5WmAu7xqtwDcjGTMz/lNdeq5eTdQug
thBF70/N9ZDDIExgzdP1+11dGcPZ8OCE5HOoR2M6RLxQeCAbXA2ptZtFULJ0kOJj0qzuiJ0UJT6i
uZWkImHg0dltIUJe9BS86Z/13oDTM4L5ZJYDKXhR1xLqm8GBw0Iy3CrHjsuNxgPVYDVoieMmRNQQ
Nr+2/IEtP7sEPfmS+VQMeud2EO0tSTG33aRUwCB7rNsaI5+pKp17KVay/URdDBis5ATSXfaBWn9E
hX1qePPK59RoVPh7GKhccf8wFnlyGhdqGMQZ2pNOZ/Jv5jX+dHZTTwDKcc+fVwCOMo1wLQYaoxr6
D1URTa4+JSi7n+K5ObSvQYz01sGMCupxWhMHS0rFwbCP1woC6W/XuoaGF/29g+Ni43RJeyK7unOf
GV6xPXsX9hHf5+cNct+wjvLrOL3k5Bn0VD3zOhAjXEdObRcFeG3gu1MwEMJycsW9WrwvMti2sWqW
s+g7tKDcoZou2efSJIVm/QlhN2U34BvhRpwN/PhGW8aMpcWCGb8phVZkCF5fRIGnsiMIdm2BTO1d
3UeMgJJBfbZHiFqSBfESnH/jJE9595bZ0nZHo0w6W+XcSnXkev1yb7uH8xbsUEu/hwNQmJLlmMvA
YPe4/R7oQXrc9CUnJp7S02QYU03PpGnQtU6tOTqG0CUYGK7t68fo3iJXi12diex9TzGQ8J8RBmI4
7F/igbH3MLWPV0TEZvzHdLxAs5IcM4+YtSwJ9HGWeHguTK3i8OyICGQHDoIgbE+XGSp6JwZuv4gN
H3AIonQ0rcuk4BN8DqYGT7gK63/7SxVjMrimUEupHo/DKufxAnXftjZ4g6rbWhvNgeeaKbV/oNxd
GgiR4IxWlnc55nZwT7cPZIgEj4ckkCh3ICfaS/LUgVI/VS71OUKQQHzYQRa/Ry0xk9IKiWRBJu7R
n1YhFYfZVmjH3z+0bgczqNWKuyxSf/NhowFrwg09OwFfaWyaRgdm1RV9Y+DBtBCc3WQX7i2irx6H
UI9AYg5DhSPlQ45V9ta+r20kcAimqqnW3SKVQLMJxm+2vaI/RQSVsJ6yyNqqs/50xXwEYGvkCoIJ
YW8a60G2zFOyL76ybzgxztNNxpPS70Z8THnTMmEtI98Rni9QUryCv/HwUFNTIv+uZcLyCFkgRqKy
XDsUv0lgjhiNfBPYQ9rBHgzopYeIhThwraFctDlPbVggVUnPjZa6229Me6ukZpiAKxa2Aweboazw
K5FWZCHNLR/rENVj2EFsVcAXptKtbOfFtIo6ZavWflFapX3LbM+8yECmvuLd9zlVhv/8RA6dodhW
OlaqELHvFY7oZgEA4HjPXxsL4gr5rHwgW8nh9F819vpD5eM9AmGimgYmTJ5uEUbJ9OcYeYO3Wtdq
H5lxu4EoQyiGAX/Ye6fnC0/HXwN2R3VPr001b+EwaXkifuLPM1Xw3Ohjw13T2X0+QI/aDKv3Eslf
GrXMntrjzZnelofKguLigcFwiPrdjTr8M7+d3Yhwk0WsJJ7WyqW25dOYWDnc/nLs6t7GxdtLxhip
CVxqRSRd3YamyyFQ9kHEzdT2GYOxMULAZ5aHCnwQ8nshYlM9wXGZqO/GA3hL7g/lThh4q//Cwu+/
8B+ZddHlt32Iy8lTRY0p9L7UYKWgLE+m3oITK0zziFXSat8+bcxW3M78pCj1RAksOpjQV6vM+Ic8
Ngy4OzktsvAnTfuUH46K25A5DXurGZa4ZOtsK7s7DgyHBD71j/9zdOFks1QzybaVx5mXXilvowC2
H3EBSnYEGVh7LvyqkZ3iIdPxV/f9qaa8MBBnTN63A/vQdUMppSCqhx+SDNpsjnndLrfYcnXQ8C78
gQ4Pwij49GsACZFia0X0ucSi1n5CaKNr7xjyCNun63XN6Gyx+uldBewLwpq5mGMP9acTCaB6NdGY
rYvdjZbzfmukw8PwEV+IL/DbaOt7YTAyGMQ8kW9g5vd98P+u9G+7MN3XOnhgENDxF/r7kXqKRFI4
Qzf/Sxa84F/bEjNcNS/8A/DgOh2t6IPNl3cszkHUtHtn3EoqOYWJMJQoZfJXSD6oQT3foUeyekz3
gMjE4ZRxUkOW3TRIohc/GhFkJyr3zS0BnVbPYtCRXDYoOAYFM3kYUeEh7ugNFDhRqlmAdGiHFQDX
1CHqgk7rkQt/umNGbBFggdRg0eZa04XWLVyX0j77q/Py6cTlbYsOneLcL7ACF2Os3pL2VXOm7wn2
AvzvOkOKyoPFJ6FfUFOsGCagBXbgm+2vWBSz068Up4OAXe11QgClkxy65zFI4q7BHI9xaZU0RI41
H/M1QWwpklp6nVuo6SjlSisvuTNw3n+jXlq6E8WK14yI8i7E0swj4pidfkbUta3AA/msdf+ttsGU
QyC1C6LkzGEEgriXEtoEGFBlWburpkEaaMPMa/lpPS4EHtSm3ar4aCaHJPAMMR5tAdcXNhUErZxT
y7VkyzxyuIPqoAElUTpgl5o+lrmrw4c4Dgbh4NyTXJVK9YoJbdeBgRgD+WmumHsPg18jE+fKRQJG
820N2jw/T6rDukj/BwoDNfflbguCwHqN3q9RwcHtHwQR2jhVizNiOuustosHoWGiN0PCatqD8XLn
WNcpsSNcOpNuYYK60sbnP5RoQg1umD9pywlB65+qnShKcVFlSJ0ZgyGGPpSSUGGYE7Xs4FXiNgGY
fdlxHSUAtqjE1ZCXf/UACJWkkmEXvjBwz/I9Wb8KCglu8rj9kHds8lA98ssOoGJIiRdcnDxYawSr
y6a5/i0enIxGPf6s3hRZhA4YfUX4m5RSNOzwbualDircasy+1+Cj76CHZtXz90okPQakCebsnl2n
ar6IjiCNXjiG514ZEH+vj26eBa+Tr1cQuLc8huQK7ZHCdhtH8kws02aoqMxVifWVRH1Sp9v49zhm
1fEgSkOWhK8sK2YOCdGpga6OYxJXXNWqZDpBuV/DZsufz7QFZn6M6abhT2/HZvgEpWb13IMNigE7
MtMlSznMbg75sJ/MjAobtBF8LSifTF8sHiyMqo055h68kzwryfymy6MbvhJabNhkvSB47X0Uq0aI
yEUgZIozVHQZbKRNJ0RVY8aw5A/wnOOzb/8e9VR+GB7k1DMkjnA1cfkAJne0d+iIBKudQgI6njX2
Wzd8SSsxaWygLnqxlLI38RkWd6UieVPmbNkoo3wgfBkxmgH7ARV4Dr7R0FDtM7blVFGnlw6r7qsR
23Ao1LdaT0u/nrQSShQVKkepLCW2UyVNGD21vU7KmH4VNApPVcrUAf1t2A6UfQmQvWBXClt/Ej+v
enPX8krMgbm6RThe8x7zL0ZeJWtkhq6uWlaKRgp9jhCllfGu0KTblXXTMMaxDSNpmZ+2ucGLug5a
UDcQ3sMCl4GmNG5guo+U1vbIAyOlm1emjN1WUhOrXT0wNBTFuE47YyvaSoPazo9Aggiq6OBPWRaF
yWAyObGAiDqykudf58HrqYfqxIfl0LO1TzJ/UA80r7f0rRCD4fShEkSQ1fC6XbQLNyNU1ilaQrWB
s7FbUXqG6TB+DRYqoVVzzIEz7fnRRxCg4kcswXzyzl+VRkm+5a82RT4Ut6PXv6U3VjyZKDbo6dDY
ESQ9JpWP9Ua/cuNTfoRdR/z2YShvD0AnMxFBNhkYJCPXCSbmsIWKX2PKpK3mdvtRY4ierOYDjeIa
iBI4n4y8cxT7ev6M1l4fsL/8O+85inajjrUnyV9jbaHkn7nGBlAWOfQ3+JNlgvc34dMqgNuKVkCC
rvKQ6K+HQeGvMJpygsZ/rJTFrjhEFsWi2UWOlKwipWFmebGbsluNPEMRIn8IvZUeVvWOSX6FGQzY
WQq8956a1H3IknGnP39QT54y0lolc5n8CfdxiG67YqL7VEVb4LfYfW34QCiurO4zEF93MpE5s9uV
TYjm8NCaepk2TahZEDnvGvn63ZPZwBACUFyAs03QT46xtt9h6SaKrIpO1KCC9EgaS85lsIJBahXN
88vAVmYmG/uHkXCjSAVYD9A6Mh84WoLidauPq2B3K/D8bF1TOxxNPiSwFq9pU2gYB3lAoO2q+8Qp
23FAoCI3+aFwNSTyGGQvQqha/rENAc0g8JHoBfbI+nDnhZx8ArBh8jscKr3s0HX212r5aMBBlfjC
YGDmqBGeWw9IjwLb/B0I+0w5kUAzICeGzZcNq6IvHmqyoi3FT/OSmew+bd9ExtgSFN5JYH0Yf9M+
jzJG0S0sP8wnENudeyrxkbFi+kW8DcBnBtos7mrLjQPyWHgPXoNFXUg75bT9fXA7+xu9nyt4BAdU
FHJXb9QbyCLMuRTSEg8EZLX3fzi4Z/rjIiRAEF2DVT3I8PF7Nk04mcbkd/j6QI7RYapyDHc5zIrd
R5Ik8f7q3bzE/Uks3vL8/MvAsodftvJ7C3GnD0JpJTsfXUMqI96AHAD8y95JQvhLl9JMIckkbyAw
WziwWmdcF+g3b/XinXkUC6ST2AmRgFxgfy8mmtEt+gSMeOnWweH8D8WX6DNX2xBKhTMhabbxO1kx
RntM2tPq4RfRxfYKHC4d/GqjhFCfrqBd7s+qg6SRmKYuQHk0jNuRSGnyYsWpdgolOgzJDKcgW/Q8
7WkQ5j3ryrkw4Ne/oSNQd9UYNQ2WMd9E/MX/6rDJOR7WMClHG55fq2kxnJCUNZTsSe5IcLl88FQm
dNU+df3EREaIaj8BomulB83zueWefQmuGWiMn/N9KG2E9nfiNErXdFLuDwv6g+lUDEoWYOpvU91p
v194GXrcPpzSdgv5/jdbWxsikpan1lNQESMRulQClQMFr4pqpMqZcJFolgqnrqJnfhM8wx2NdJjR
QV4ASNpq14j5NsOP7eDr2FK7dNMDTC4UYg4gC90XW2IRA82NsxiE/DqUl8esrN9nCHGsBbsDdptx
uoUQurV8tolPaLuZO0VpgAJ9Q6QUH7Vv5/blXook+dLM474RAo2GaXMTawCiBTGK2EU0MwUAFlLU
vK8Wc44Qq9wuIBZZ2Ge4aBEoTNIgohC7bbcTBwuOslG6aYG6/pYCh1Zf3wNiuZkndnOsb+WRz0Cq
/wDDiHB2OOuHB3BlJTzM1RV5MA3J703+kfj/3uVclZEXOoRUI2IttfdSFRwxQr+WPcI+zzzZXdmS
LxPAUap/0da3OtmxB8/XVFzhcNnpaCDVPEIJJ9L+qL7x1pYk349vI9+QQXWbIzpmQDTvlNeRMaGB
c6Wmb6xjQxZwSmOEQhwDajBJmDHufed/2gLeJopGbSWC/7NN4BusNG3KZ8EbU+jIgvyXzcPGPkeN
dyKyCywkvpL0tIvQNcgP7tjYat4hzTGJ2IaOv90o5DidL66tF54nTXTREZe2CZ80tMbzliBvg0Jq
MqIY1t7WlDEj5vb/YUKSHzwtWDXWWp7TWQzpdxZ+OALkCZM15D1VG8ajUNilaOIbL5QHC4HjaUn/
DKk+a5JU/NJgtGftEl53BupLJUxNEzRehL2OX5mcJ3lNWdcYObF1G6RHlWFZyd9lW30MZSmza0MW
anIBmeit23XWEqZonR/zoqBkczfNjpCeR51YJMqF19fIwnPvSh+1+YAFgXvsMqZAeLtYj0/WgyY8
OSvR7FmTPFIc7u5bgtbe/16aCwQGfC5JZcx/1m1IbkFl65w+PJHWcHiNf+YsxMhlVO5xNHwSTT0z
M498laTptGTRgVkPMh2RsSS4R0e2AbvBWSnNx+9UpMy6mnR2t9rbyfwWPkIYoy6HU6XbII7yypAi
pkrf/85Q9U3V1FU1X74ob5Ss94BBYCD7pPvYFk7u08i6lKnz8k1iERz5b/Y4ea1Hg3kIBWTqz5mX
bGLz35mIjXEsPdKumN4u4v44SZm9vs9sWH71UIzNN6o8s8PvfqyxpNs/wo9lhACsonpj/csbh7I+
Md/M3WDMsPKYAoMTl+jQ0PRqCYGzWunwgED0nai2AusAkuu3XI7rAklSJVeMJAdTAWH4beR3+5Kj
jM/yt7tPPlfp8CGSAw8hE589yKLe66lOjgempFK1GSxkatNk+nnW9Udyx4a3tUPn+akSxADVvFje
fkd7eI6oWmccwjT5nFOOu7F/z7aq9QWsSJCc+QuS0RrzWTgEvlEdw9V+QHNtS11uFvlpsYxKKegT
H6vlsX/nWaopxZWmLO4qQ2w5OtEohOk/M7QflR5uA16C9OgQyPmglwEF9xvucPd66oU5kg/DFz6i
qarbqkUvL1G51ScrsblyUjJCPjhPJGxiDnDVpK2C8h9fKfIoo3HC081HMsSTDj7VLI0sJtOEBfL9
maMhEN+gw+yTatr8VxyjA/hd1779c36nzh7WKj/bqCAlimFsexQlYT3RvXl+6phSxtpGQBzaInWQ
nLEKmKwyrBfOTSzcKX0h3Oa02ra1JXPSbRVLaoLMpYzaaYfkuPEvbQmQqxKYrPe31UQBcB9VX18d
nk4Rw43qonNfMNFQON4AyflWiu8mQX2QCo/YC5Exuo0O92BcfCC3bSWSwzmsDyC2BRdsBN/4VvKS
RqpwLDTdkHvLw0AXN4U+Qhn7VrzzbLzmnokceHph8zZKprYgUrct5+04auzfnrlT3tSn8jhyR0O2
T1JI8lfzNbzChIVFDR3hx7/zYBIp6ds/CQ0mno11dBo+Hjh174Y7WQzBWgFzIKiMhOHtgcBlcIjr
0JOASqa5Hw2Q6usGfR876n8bAa1U+OFUYcruXiqvs64BIO+9sACN9l/JfGEz1Cl5/eK6uG5Rvd3a
V/fofoe65FTnTIq0hlYCmz8HdzK8njnFOASiRS7yVjXFJ6vme+W5RUDgG99Ge2LoK4zFnA5gEUFo
xd9OuWqdCPpXTXAksHsxwtOJQWC73HIIPqBfDZysDxRDYUpY7ggwwyteDnUpWp5zL62HniREtItL
MyE0jBJVHu1F5lW7ez4k9EOx+XpYrO1QEi2HGmELhp6/YzrizHUQxlrBQ+gz1waja1AHCsqCqOxr
XPAuwZNhWcpdR6nNglaNLvTa7ahIaqbO0FjH46t67gtefrHZ1O+PgCqMmDLr3fr6LS+dznN3RM1e
nl4OUK3TwQZKXb1kv8khdXrI586LcuhSBfrBNs9agJdDfJfMfPD5MWsv0sHjredoUmztTwtTrnJY
Nif/lUwH9etQM6Fjg+FLJURrkIiOuMPVfwv+0S162yjycxvj12n0tOhVKrzwHk9WJXTUJGc1MnL+
+1lndAxt05J7fMf6s6LIKxUwybcx5sIUQUMKEuuC9qSmt+q/rM2jBDDYrnU0praHKwhJYhTSd/0G
YmxEv4soiyUTc+2U4BJeTt7qpqxLmi6uSnGDLu3D66djvncZ9JbIqtFzQhuqihELr+21B7b+4YIc
tfogyH5t6ira7EYYa3A5pxHP4b3NE0qqQRIwgK4CyzhbXh00hD1cZItnim5duUYLf0SaxunWH7BR
dGxe8mqUAOZZqsCa3Qt1yXB+0HxyK20BHRNPlVJFmhosSf/tPv9avzk+Bx+lMrQHjCHQIJOak4lH
1oZFxd633lVWWrUcAZ6A1+rv+0PIcevmKIByGOmeOUpPU1P879QD+BQAvhNvfTaqEdSkJqZPtXgw
qCX3Z62/W/9n4tgWl5fuCdyJMkfGyuIxgU70kgDYIOCHtEJj0hSi9+uPOiUeLvTEa5CXJNNrWF3s
m+GMX7je2j31om3y6q80RRIV8QRBxeq0sbYiX56Gisy2MmBuYCEBrZaTWe1ck5or/Kg2W9Uoojta
lHzTfIJHRGQ9jhfKzPPP3ly6uuKEYAealT/s7/abTl7atlS5D+OwWmWlPc4o3AQZpsBVq7F6WPw3
SNrgwv7qmky/CWe5r5OhwWaQtdN2/pYRWoqtMRcNcdI9BDVj+5RI0ulLnHO9PHe1QMoY5RWyzBAh
c9z0g5sFvtaS4OJ1GWC7h8FDdn9S+8qf5XjD1060lbYbid77Cisc1GHA78+oKiVyCb79amKG3Nwo
dlpKF45f/qoDz8b8n9UIT0gQSBf4hMSlG2NyHT0Gv1ld80B9h/eTEqcajABS0AhuqIabwfR5hh/z
BnF9+juj7ZqyL/1HW7uqMbCLgHwGRLeTgLB9q17D96i7MtFsr8ws6USj2dND9Nf6hMGZwtP2sow1
AzUlhy0T3a2x3R+SWvquvnFp1I6iNpzFRDycrc81m1y7oXArPIn3wZHS3nQu4TMoTiVOf4jqTNl/
QUdbzQbvlE9WC5kXxybqd/u4Avw8x3HHC7OCn8edijDfD7gxpdFYAzXouIND6tc3Pvbnjgn8y+DY
DqifbtHxHqFlWOcRR2RTPv17quKF86et9zDO7v2vcfT1WA6G9JgZHbjTrPzdLGVPV0/RT0ueIKbP
wTM2NbAc8BK9wDBs4SshvMo992++luAJDpo7jAKTnh5kyFTx/GT7HkYmTxEILiauO+j2UHXm2mJz
yx7wru37APc6dCp7lTX96QxrywCFb7HnsGz51qepDAh32HbJmPkT1xH0IuHkEAtgw2wLAXQER7PS
D5NUTF+W0HFeKI4nlXUFkn+Jf3NzGhXy4YScbju6CU+X0TncnBJ7elB8E8qAkXcm5SG72/DqtqVU
vcx9zz/N0b8hgzghbwpksI9NKdDcdgnGGgZM9Yn7cDpxc+GTaW+qfxLzqSoKvbvFlcC2kr/EsowP
jJYchZZ29icNXfrkqcZ33EWLwDHgrzSB8UnRWvEwQkjfDWPafj7HXNxzhQN2uye0EtvZekPIAY9J
6JyPPVffCp41BWeGcFsv2hgLWikJ6fdhaIO1/vzari2Fi7ZCOwyNJYjZ/b+7dYJF7IGMco7Y6Mxy
lyKJ7uNKtSazgkT7dl2HsIdeiIfEJrZacVhB+iNoRtyKnBGLiIz59eeyQ1WMnGeKtkL1OqhXB23u
hwLnpo6OKEcXcwtp2sOF3WuqDWxMDSTGmZcFoD5D3NsgYPBIWqrndxzcET6zb82K5OC45BvACDIJ
M+gyPx5fG0j05XFPRFN0D0vwf4ePWfyE9uEOugQeztlssnsbUC7m3BvzE5Y8NfMRlcORq2I5ELlp
55ektuVNd3Vk1ds75AmD1oQtIttaEtgp6vaeh5T1IxLhAUHyLC+rGHhTIqurDtm/sr24FIktdBhg
3sq7ullCDF3MKMUtiCU4Dg1IBWUL6PuUgAvpPQNturvuQn1lKt13OCWfQG3mMpqoT5HoN5P6GCu5
UczgC/4yJtADKg0LDec0YUYUKMu/fKqp/vG9aUKSZOFLjxqC9dwsfTTwBwTGY/sjXPh7uuj7wxWn
oQc8yeMilkQ+tJw9xg9TTg1OZAjHDRf+RojS03YeTj02Vl01WE508SYkXqxxEphLZ3oyW5f5cN2T
VIVjgcwCFc68Z+RuSCF4SFfLiBYb7Y/W/d8XjyqQ8rRAsIMTZJzjvgDlnhWnCPSmlGiMOotkiAWs
bl5Qhyw7fYNhHcyO0+DF/MQXGVGlkgDkeyAb1ebmshMcP1JdXAZ5AHKm7I1dkpc6a9B2zPAMZ55i
99NGxThMKET3b7CL2EDIxvkl63+3Wx6GeBDO5sa5JIr0+sCD51o2gTVJXplQv/pqp+HfKc0PcS1I
3WPhSKu9Dv10ddE+ag6EjhtZpSdYgmwHC5TrgjvrmJ0XxvRUnwZP4ww2l9ouxWEH3tlktk9JV5EC
5hFdiWRsBDBcyRXy3WWjzCFXinqF8u9/koMOTfEAcIHndqfsX8d8ESL4Kuyw1llYkielDQ8EuMns
qdBSHwPvosmN77EPS9ZL6LMOzKgLqtnNL4XEVGuxSmwVN1plICRa/zC2sIwbVspensMOJKRb9c8f
DZRQNI7Qoge3Omv4cXtMonflHmG+0QUy4ekTJo3h949YIXvZQ47p6YdjAelyKMsoKtZsVtrDDry2
hUCvJ7ft3IlAhHP+UNtnCUPlYKAOHr5ERDdLNwRCGrb69UxgSOdfrBxxOUYM5im9kjiSLEC2jIg6
NSWQlleSk2CmmqpvTAXCzg35E+XQ5DLN4FcRunTCjzg3fh875Z6RBXWsUgi1YAWvG8c3JOw6sNi8
urw6FVhxPToqWpW/EkyGm3gw7g3M+ZhpCzzkzmEd+Zb2+0+h03dddrm/iP+GQhAp4SXyCQQkZgTO
Wat38R+ACaLb8trR1oYkFuxCeRvvQV4rlMJeHSaVwH8O34+96+wMtj0KZmp/zGj8jjHSbl0sLvWI
HaE5tigCPFytSOuB1jOnWJAswTtbqdquOHzElemlQ57IBM2Kz3JkJFIO4NEMPUf+rTzCdzlCBByx
R7zRc9WrBDEaCmTfEe15hl+pScajlLDf39RQG2FrFaJALjguubDwnk+RlOj4La/dCtX7h4TN+Gmr
7LS5dtXycNIyA7j5gUwZ8TrRgVPhbnW/JEak0TpegkPffkS/3ORgOQP1bgpAJjVDrL+w9tdO4DK9
D94DgXE+apQuD7QQHjmf3c13sXfA2TWAbrpMNXoYzDfrDCWALdPKHD464z64pt3503DlHscPLWxp
mXAHo7vBmXQptgUapYxvjmOtM7oNEdaX1jboJxPwBqqvUH+VYof+SRF2zMo1RjxCjsWL0ByFx6T3
zxs/OZA+NLatyxqCMMhfT3AgDQc2CVsfldUfVJXyXo97e7vcHrK/wUbbnRexYLfMVkA+SmqszfCE
l97HIVxRGh092X0HLCrfuE6hrDVbH3ZfJtAqdzJwrAOda0UQBvG8rq1uX8S0wJCEld36PVtBbuVK
S1jHEEApV7u4rHYK2cQgSXu8EE1p/MrhKq/H4PlwacjsbXliYkLVYYwXY0hsCbU0rHgf4EMp9e02
djXhc5LDIwu2X3GuIhPu0szAid6GVF9wrYZ7KApLq3iUX+xp6YcdbpXd0Jp6DqUPML3K/A3lpRYo
u7fZ31oUVTtcFxLHNa28J/1n1chPiSIWOMyOD065yq/gYwCgt1S8NMKJL4b5zwkgD8mHsrN+a85f
zyFZH97cU+L4uTxpB4VWYaZsTtHA9EoxJNcptyvbvFUzVQRxow1dynZuwtoYO8j1dOrdOnk6f7y8
6VT+m7NTEcbtLYFGr1YUhxd3kXP71k8VNehGeYyyGcSkacxTXyTsvQqV8q5bhoYwUM0tdL41mXmQ
XXcUzCobe0Uay1X7OTNOUSxP5kZCCt0RvSZCapDXzFKJ4dwviQpnBo1cKCwudeG72WYTjRwUB+AV
UhHnnUiz7SwXDyG4aw4z9XzxllATHo5uBO9GAyTe4liZWK00Zq8TmU7T6Lhd4NcxFl763NqXjGH/
1ud4Fb9qEoJ9P0aIKayPUoktlidxRiZfi4DSZvok8BF34iXYoWtv/DfiXW4gvz3Bjp70YmvmxSVA
IRjO6CUSmxQPDAiriMLCXWM6Haxoqh69u6nEN8pLtTcIL1kVzcrZJWXrTVoFjzV3M5bxKE1TtTci
WZjHpmkcGhYk3bY5SAHILwpJmb/C+4MxjnY5WVPJD6mmH3SCr3EOSVKT0RcmMlGUR3Fcl49RLVo0
TuXbfHp7VRaNFrYYtm8feSB/Y6/TscZzAz/ZQxMCECuVJ0cO06RJS8v5DUtxwIC9YiGj/ZkvW7pU
tkrbZhaxIF1YyvL1C3ZRP8Vve+ugOhVhEFsuwNkm5cWSpaBd/PO4ezHBgDsRDIrif/TFXQ/2YCoz
7w3b92kAekWtzV8eK8kHsj5wdog0sxm/j1hguqMsZxPmDOr8um80nFUrVTc8SsD3FV9poRdZ95QF
FdKvylqGT/93elLe7OonKr3dgKwgqI4cyBbtxT584b3UTTiZO06xiQRAQmw1+qRibuYaDz5VZWvI
o5x8Ojt+143afkSM2y7SFjVs5StRyBe3Z4frRPfL80qMn6jVoya89lighniisaF7rN1mUgNk/4Pn
gQ+jQyWfEBTaOMbXd39tB1e4i5nCV1FY+Fk+RTDXzvAWgrfkMLQI15H7TqcU5uQ4eCTkFiqowmgX
ZuRWMLYSAVM5i3mGLlJCYB9jsrfonXG+XMfLmriYrIeB703a/yPEZAY9fpgdtsB6CDNMnZ3u30WL
V/QBGnrH0GQj6cwV3lViFLFfIGpTosgVg5s9CS9BZbXJjp3dskp1tfwFK/2eN55K88OFFcxDV0PO
IF2BOcln5UXNFHSZ/sqjyL0/FVc54Wl0cVu+46ChomcBIKtk5paRDK6dqAzNGUZ6dvrmKYBAGv35
bF9U5Ko9gyD9ombu2/K82WwFOh83HU0aD/MfvNnqKpDAZHhMWSRUOrk+CHOz2NHRNQ5HtpPML+p6
ncR/9DkWtoDYOEjiv9AIK3tbc03/23mKh5dkp46vu35bOgIey7K7fkro0lo1S61KV8jODfkTkdHp
k0eDuYZoEgBvPTb4wAypqvVs5oiLh7PlzR13FzintimmM9ohHoHlx6P2ElzlR2GUfWkgPNCPkXRf
mFAuRj9oeEhDn0qSIwlfDK+IjNtSAnDkFF/ziiOS8X7yLVLxkYu9tEd0N9mJ3dMARfUn/et4b/S9
qNzXoWNgOJU0JEfk1SAUe8o7B39xnoE2sGZAxgXhOJe9fyt19z8ZrDCezFxraPQTJyVHIs+xKsVn
xSbouS+v0PjWfMIMGrK1nkOtTUDAWF+6zDlKvO3c801IzimyRr04TOLYYNFJvC5pLURSb73ssT0b
UdVE5swhohyGPP713yMXEXpqmfw1R/DblbFLVgFUxTthZCE1s9vRbTDUPJnrZbOHZROmeub9IDkI
4KrSBjh57yDqVpocDtVSx+K+PHQqUYbGD3ZHENBo2yEVGCz79vIhWCQYQisa1j82VyNxYbH9SjRE
e23du8vCe4I/r0lGva/CGrfexAeZf8bTiUVY2Hesp0jk+nZgy9y/DqeEtTtnn/A0V4KuuQawojrU
4rCwzySgghb4VkJftYIXBLff64LN2uveLgxEog9j670Sb9BwWWbxHLqr8P/EmQs3Nw4NSRCRFMq0
yrPT8VqOrP8ctfb5b4b5tj+2L0AENP9PtuzGZ2MwoxVNcqnQivC4+VrT+VG0lbOhQTsWuwXtu+/5
pBH0GjGz5fHFIuf8cRVouAJP3VboQySA1D3biXBYPVxwvdQV3ml2HCVMAmHYZDF1BUKMG7B7YVCH
fDJYXLBStz2Td5dMgP3TZ168V9rAnAYkFFW09XNQTFEHPBKtNzqys/C5+BqwC03XZdVHnQtxJEnN
3GVPnTPkvvH7tv+xhMPnBQiW1GvhCTwDimdtpMXuoreeKxB+paW+2fFyJVeCmI7LInvd4x6MXQ3C
otkMmyXKpbkCXwKfOpKEcMZqdjBbYFK49E8qbt5OhsdChEQSKW1Inruq0bjY873YiBFLhku2clhb
/egLJSXow0T6frsZ/n+5KNaLhi9dOyHSyuZjO6R6NmorucqdPYqhfK2hEndaWVLLkMQDBDizSWz1
H5r6IgYoQRoF2/k6ikoiqCkwQzLQPFpQ6z7uePl+rB7U/WxScrhszjGYr85DQfgjChPsqS8Zgvpz
OzEwudUdbgTV/+1Vb2Y3jWWplXzCfpPixPG89q4m4HkyOS4Rn2XZP/O7RXQsgjaTmbeuTVbomIb+
qloaDOb3Ti0kWHTkNRrUiY4aw4XxBEqrhsNc7C4mYhhWGXy1TO3t7VSWJV7noefW+rtus9a8LYsU
fhFvCIlAQbgNNwK9vwFFh3Y3+G8mCW2t0l3/utD/Lkc1MRWZNV+Ws0y/bq9jvAv+2eq/4NT8jOpo
Uu6Irt1QjfEI1iUP9+gRSSeCx9PvCoUy4dmcCJpsAgI9smyxWVlH38bFJarrv147H46yDcXFqpG1
AQg3EVnYB060wB3QFS0cBZo7e+YuArv0XRm4BWs3sT7Iux2VqKVfRbSyhTeJ/Y2lPf+LvEsB6UCJ
dkONvde/ISh1Ek4C+F1eKCfLQmdyMugtzUr27wJ7EIVEVSHcQKB9ntlM0IaK9EbvtdPZErRgq4ef
IW1y/WmdAJaN5qSGqOBEgNiSUyUZ1wSa6s92a1b46aGdF4sq2qMfnXYmqxp9ULlV1khs6SvfxYBc
6O+3A7lm5rEZ5H1pj6V6te3GaFOibdnB03W/eWzi7pyDz8pXQlwk2gh4GiOTYc7wDWYvZz5loKkN
/fR5J/8UIUtP/5SV9tjwFDSbuAELoE8m2eoMoyr8TsBtmkRHkvHRH2ChcVZvsi0cvC2mz2McNtYE
3jD/otYPwbuznnTY1X+O/11mrRtaKY09SxxHq9f/VsVYV0aWXhKiNKSx0TLJ2hj3REFN/+ei/Ula
tf8FVF7/7lAAde68pETQKo3I7eSO/q46MYNYW89SpGXXtih8mcaZQ24yO8WB6/IYN+bqDZFvXcW9
8PdsENE78FaIvnwh5ookNVTGmrOjTSeBIoOp3ZYRTg4OOElmrs0ruFkFDhWnZ61XHIW178RRtAam
8VibW3Xc2qlffBBT0Z5ipLPtGBlqK+D0jyfE4nyLN6xqrxVdREC4+hXHa2HnK3HzXC7t4/O+UIMJ
U0hxYcMZL+2fzHp1VUYFvOnHYKXwFIXfHldHdMQoNC3ooXovkcIjrcikRbh5Rz6mG4iFZ+ItOiY/
AZEtdfpKworo8k0R4Wni0UPbsc2CXYwp1z9teKnHG6nbNIKZP+5t18idE04c86Ent6gsCZT7bCUO
tFsh4XsIRHbNjLx4wwjtB+dRVg4iLr87hCF0PHXrRrykp8S4PH2udVkq59MpE9gCQaakOdgBvv22
Sz2NZPDCILTEqffxLqiENBpTwk8usys8v7w57Xh+vga5dFJek15SiYwfmcEQJK7Uj6uZ1T68VexN
Y130Z4H1c772iLBLK8gwDz3qcxyR3n0JC+F0y701y6Y3BImicTD2vVnIaFyQ80Ttg0/4gEZiNqg0
BAw63icTbzUG6pbfsMqL+kYxsw1WJyQfEwqmMc6LPAnzutsGVoub3Cty64R6VVYXOdQktIZHO7Cd
SVc04K5PUh68F+1HbY/EKcppJnyzinZysiNV+STcDhBJB/BvoLsEib9kEWXYkudNeYpFXtlfquD4
y4DfLxwXGXTnQUiZMGFcB3flpyf2SXXOsAAdMMsm+9lJ4l9CaeWnT03d7nQwc7l4EhsLD18VOXFV
Ad+ZbpU2Y6iSv8+gEkqYM1n5RQSlQxUCJOd/Hgkcxmp3AySnmJQCIBSebfueUfGmsztawCdsPGr9
s9/CI2PSgLTBexzpwl2mjDoEoAofQ5POb1nlx7+9Rq4q5baAQhyRiqqE4nfZ6tI4LvFrUy5FfA9n
QE7AkOy5lQPbMTYs1lrhZ+HvSnbFEhUPX82yu6KQJuD2+UT8k0bSFNp3Z4qwQrqnvkz1rQLBrAqm
QYmf5tGHXYVAjlXuF6zxdGfFyaCS6l8C2HCdwTYOOTSbi4FwYEtbMHxB0TdT6fLEVK2ChpU+wrIO
xeSSoWimNZx56ld1eL+dWbrhj8czyl42D41mcuNiy34oNGbfpg/Z/JzbRf1oWT0BWtOv4F6I+dtE
qu1Yl9jDVw8hWAU/XPUJ2J/ZvKy6yR3/Fgap41O5G0TRW8zkdEN88IG2x3M1EZ5U08+XSSTUEupB
+aKLtIaZdk1mp5xMErGlkUGQSBiQ2VSlsNQ/UK8qhqRfQaXcvZLDzFbSe3QjAYiLOirBssXP84h1
jexmrfwENBCImDZgqyUp7BZjc809s65G7HCM/UHrLPo6b3L6hnpGpQ0yCBdCI02yLlmk1uRCbM/4
0ZP9FzEQa7ZmPrRBpCRJSL1njzMSyX8N6etlsq0o9Ve3F7KtFrFx/XJhYlMVpX2LBGcK+1Cma7wc
vJKhNghxHY5via3d8f/jH1AkJ3XVncKMaK5R8+7IIeI360azGbh4Xdetiwvnuxm8i95MalriIYhY
/MBBreoHdPt6RbEIIqYxPVRQDZVSSunbxz33i8tN00JJn5ea1jdyckDs/vjaJsExPFmB/Xh46S7w
ls2VyZ0WbfR0yiACr02EzshEWBEt4FjmYa8fenO9gF90d3Wf5ETbc4WZuxzAJ2G3sIhg3L4by7sf
chje4Zzhl0vQ0OnWSgnNw0mm44eVJELXDIbI9ngjak+XPhJ4PZi/1j+OcVVutK+xeg0KgCxhOaxI
MGHzUcrNo3iioLJhz9C49cod5xJRIKHY39m0xxUyu7iN2xsVHBiY6Qex7N57OTBCx+sdWCsadX9P
TiJX903e0aq6T5luWOKok8R8ZvAUvmBQv2CLO5Rm9wdd0wGgYLnu2BBbxSgksD7dWPQUkcy0GRAw
xcR6wxf4/IsTAvYltq0x/DIXEVeKz/q4L1lR1zgIb6fypGPebFiQd9/HNhm/QkHKDyn7spcmYBkZ
F88V6tsa0YV3tOjrIbudwg/rTUjaxWJYcO/s+KT91JmhYoXI8Vc3xf6ZYP71MFR9pkJKBmFnPRpe
sDycqsatJT1fp0DGecMdo/3WgsqRReOsBJXZNAUUzWNPFt7bVDt574SSNAiq+NFEPdRNNRYtszYc
/960LjWMb2VvqaXFa4Z1qBarjds0kKcIC5czNRuLfHickRxhJZz9DyPB5RCz1aDSHvgpR4adEye1
ncQi9gLrcYR0XCncgBofkhK63k6kPlDzqJxTWTXwvnLEYnFSZOjfToh+V20t/OmGsnAIC2uE+hD5
6JmoIsB6L8Jlqy8zuHj5hXVG8G4vwtH/vcG4O95P9RPW7k4U5crT9ADn8oAEv6L7/WVNFBOsoRVZ
QJY9UflYxmgbQtlQnK1eNSfyFwibnmd/gkIk7WNXfrLbNybzXtGFp1aPIT9cwdIwCpAjIK6UruzZ
oyD5KPe4UfHVUDVNY4/Wfn9MBnzaJOMux7QRMpdPCLOSp5Xr5npeK6WO6BvdXPOZt7WMy1nTgp/z
Cy4gVwXM1dQHoEdmKPKshp5QoXyqZmlRhSQlkFaQmg2RKR+kAz3yPoEQDYpdFfGdJXsp6UmLLcZX
MbFo58Yj1BGvE2FBuCyI9+Ffq8OAVYEZKlQuQOYvhQrGskYYQBt+mCJIuQtIZJB5Lx5TSoadCxLh
gfiYssHx4kLdaWkrPtkT/LCGDNSmS4jxUo2SU5HDEZk6NqOR8Xiqpb94AOsHVCsoXp5tb1qfT1Kc
mTm9L+jYqgaZ7CLHtYMuxcQHVwgGRxW44f2aexVAcfv3PEcq5EYekMvHQR7qtLBUtnkssyxkfSja
7166BmfXiaCe7WhzWCcrrBPa4LDFzEj18C2LmDn+FPSzAeN4vwb1znScduIwZcIlZI9F4Kk0v8qR
aEcLURnWaD90Thl/dn58Z0DeBnN5Rx/4ejudmA2CQajIhLPvPtciY01p+nH0i+JtGtzQbYYIMjQ4
LyKjbBHrsC6pu9nbFvVK43UbhiJJ16G2OyGcfPvev44DmTh1p7u5lI6ckkWqoYn+Ta0aBAzZ2/90
+QWT12vn5yEpp6mo+V6dqe+R0fHFSLDSLf/EFWi0JhE7NfaBK/8y/+6ct1+FhL4vBCCY/gzqD4HJ
5y2rrmXcPjBELjK8sSYgtDuehh+Jedlf+JWCkSqe7ipkLu0xIeij4yoKy8t9nXE0RE0vAYO2k1XY
zauYqZ2chNaPiQi+hJ6cHVJXjoUONgimtZOBu911EQ42sfPJd8in2q7+ykkssxl/WZMRPgYTRIBP
oiHvxYuNOafzcx92UeFrs4m+4VAfE9Lt9U6gJlv0iEgCG1y/JDIpIp83Hz6NxDKSmOYR5RxPj2Gs
ohrcqq+xfg8kWXMWJ/Y7ctHEt4r6m1zlABqN+Auoyft5OhbWN1lG11lS6frzio8iXLPwFrsaABW1
Rr+pYEtdQCwRAuKmsq8vJKjQg0JxhYjfZeDs010MN+oNgjNQDoWV2C+BCyLE66oDODKjHt5I+Oq1
kFma6OK1Gn6zwHT83QiooDNgAI1LgPrjTuxk6Xk2ML8r/sFLrDkSAFKVxNTa/B+ZBp17zo9oJjXR
sGItvGeuazK99F109WgxeCqyTPXBvOdVyMG/qfLc+nXDX+/bsEW0UbLST15dIj6Ark7Hhkejp2wi
UW0p+rvjJJZ58tjRNhxs++hLl2rbXXBfPKijOBK0CSANCkKJGcRXJ3gt6cvwMFAVLn6Hv1ZYT1Zi
OruBN9sRJXJAOBG4v1pKv3OYyUdl2mLmhWUdfhbwW9hzcyf+hbmGsD4PlREQamB3EemJb+QNnc7F
IPNZewyCc2Sohnwofj5lICwOsDzYWIzxbl+bz9QPaQVSWVByDoJ8aCMWxiErKdkJLlfLt3nQL6Ba
k+YzR07nBFZV/G1dmZZhOaaJ8E5VJ68dBKyRB0Cv0N1rFr/WY5hGfTlwqzSDPC86hYPW4XKEHq4n
5gfclCsbJu86LjGivzPXIYfI0zuH/0cTx4pHRYNjcJ0rGDNDHqveFZHgf/8Sc83b3COt9i+bNGEN
gtuHGhWURVRZQ8Ufq3BmTtYDR+qOmPJJ5yUSER0bhJDZ8d92Ge8KDAXwwChEVpEvcEIxlVjcYZKP
gUnpcGfVYHL49tqXv2tPpEykGYxYAzkrmvCh8yXE4FPG19uMw2IHCwpHUihm01by/ZYJq/7m+6DQ
pA+agIOWJZfBTGAxnus0JQhuimIT5Kk5xtSWHywfOkceFXdyuHTA8gEWKrpyyCjhMz3bOhqOrNnP
9xGQXCvAZxfCgwgSn/yrlKeRmUr36zWkLUCIGy1K6CJJ6/Rp00RV1bU3BNLJOwLWxCYTayhL3/5p
nVpbtcKf8SGdRFwNrQSvmRRxyUc7k+nzLLy0Ovt1MZrTGEYCA9NTlYQ2pCnBk9KM0c31sSuG/hLy
H9zOCTHztbeQ6ntOhYEg0PZhjCiJCqKQAXwZoJFa8xFKP1aqzjaNlVWeo7EhLpEg33lnOla7wA43
9VAcqrxezQ5WAMHdmNBoQBNsdjemUQs6DOSy+qlHneJlXeJteEf6V3Xd8XAkB1VnmHQN/tVTBZ22
oNlkzbNHmT8sJxvQ4J4n208N39+125jed+13pe+5y1QJFIRYi55GJK6R1EYebLBQ4AhxNV0rm6VI
/zuA5qUajZ1+7UMf7ooUGhoatr5D0VrNjKf5dr9mKiE7CcDPpBjAewHRKCltGO1SJCIjhnE0cUgc
Lz019Qh/cePp5fdwsP5kFTXtexmMx0ZX4ORRnsqUWtbLFZ4o21wOwnF9yDnmX1A+LYNjNB5Me7yH
DcVDjP8e3D1eSjvVpwYUDozkEDNGWaLwj1Cz7lFNmHi4TPX8VUXtiCcjwtFmjzdDULEEY9s1X6rC
7Zimn+CII4PLnBEEDJSrr2vav5Pq2V6SooL9GwFwYkYyv8rWPhFrYYQCoYd8sUvqrNWyvO9xSjNN
X0gKzlKfvM6F9a32Y+iIGtfQnxt45GUrAPvM+kn8WpTyeS5ZUuSTKUzkjbYxNB6yPgOgtK9YeOtD
9Bq3vB5fw2qpy6xnETuMWraMejlfN2yMvIqL2+npnRi2DlhcmW9K44lA1OxPxaUzV20I4RqG9UIc
h9b865jvsfGC71qka1qMPn3WK0hVLYsrre0uuJU7OWPYsIpJeu0wMo3Tz1DNDDR5tVc0Zko+SPuJ
BxgMkdicSUaaa6ZRrbcQmYa5y5t/v6+tCq0m4qHL1sUyFA3xE4+G0pe27b2yya5SnsGN39ixhBtG
ywQ2a8nNoh7cJUygcEGbmIC4EGNZBWlTcWPTQF/FbYnYdcs1nOs75aG4fd1+FTDQGN7n0FhhyEqc
O+0LT4DON5F3MnpUhOoKueEjrsf0Q5lW9/O0Jb6fV/BiSEkC1wZ2o+qHnoummgBr7ZdFJN3HdG2L
+BOMxXLrxXai24YhbwqEiwEsrBw5B8ldaK2MLDD7QLqCEkyEc22gWzk+GMbofy6KPC5w0POsIFzb
g6oOY67EjCpCwbvPONA9YB600KIn7ZaWytWUEfRBRqar5NrlJT4Ccn+WvTolhLQI0KDzE3ulRwu/
5ffVa3FlyC9xsWA9d7bKSGjJ3apF9wzc6YwcQpgC6xEqSlG+fcQsAcnUryqTemomLS16NqIKgKkw
rpELoRnRX2VPiHUDqFC4Jez3td8aSiXFxmYDeQWPNL6kSiPBEmrKJSvfBYQMpXj3BUsz+TmKCRHN
IKd67td04dO6BsX54SktAFrDq4VLt2dBK5q60aAr9NoIXQ8s7mOXtHR2KzOdnpoFr285nru7sdxa
/do0A9XaVVAncgMF0tY+CXG2zBiSaj1vRQAkDcnkbRxaeOUSBEBwamyJ2aN1iu5PNj6aiHI19aXz
eWhMP2c0Os4B24u89q8nyPNOF1ScJiG6npE1GBhht4hpg3WASLITrR9K1dPwmRUWlMWCrBpzrQ9w
Se83dzid8T1r/Y6EkgHg7NeNkvNJEb4I0o2giRsnJ+xXFZTxO54f/lKq1NoUXOcAAWR5uFkBITWI
2YdrdH1Gng1I39J3XlCSZkB3RC8yBheAOWw9dQEHdmRXYWuhq1SMtW/cMFUjhqo0QE0E8bDWe/r8
Y1qtVa0dpbxpogROolDR8wfJm/bxRNwDke8g5AIsNGnMBOJsQxqya+tbXZZmgpf4XpQtISRNM0sl
o/Y7ByL4XMnCcK4C6KdJHV8ZRaUlB/8vQxju4i1bz+iY27VALLyDzyosFedFl5zvj9kWAeC0E9B2
jKzirItKb3EhMMFTD7KFzRyoXqomsL3FFmchrMaEc5LTNWOm1MD5dRkvOt2yX1+mQQpJjCLd0dka
JsFrCsZFrELtDfD73t2/BqDvH46GS2JmF7WuETJL2QzTxtXscEx5Vp01xWNbf+d2Yey7aYckexpL
wR/3c7zaoJnIr75KaREzIhyZaezPzca6uJ+13RBsJPzybToXVh0GaGorN47KzEJD/OqGqqpECa/7
PXKzwXkcx5FEhaOqhZwRLhOtbxw/LNwauRh0LQL/u/pkup0M0XI/OHINb5/cugKcSpYHIrNv8KCl
zceMyvZOOc4MglNDvZYTRez8Hk/E1yns5KOJy/CK1MaxrcYOEY77L6PeB/cRPFb5m5QYQ0ImiXAs
q4UWkQwCY3aMQHdc6RRN0L0B51vhM/1Ga3ULlntabLg8zwh/fgSFQHt37LbBry99TmAY+rVsSM9E
qTZ28sNM4KIX1V6u6rCVV5i8yjzZjh/GGFbavJGSgz3RXC6l/inNPrlMeGcJvuaXTc0YnnAMmWNd
7HtvVbALLn4tj6naPQI/mNH9HBRxvDfiuL8I2r6khWhCP06N/2qhWnZHuUzDJlsVw+lriw9R8eZF
l7P4oDubNYhl1cLMXozkUpGe6aUrBeWCoJI6APDlLT/3356iDGy4NW1xR7wQzJedsl1BBkJ4mIUj
eV1jckvAI/O8nmcbi/2ncZSzCTOIUbI9NGvS65hzVh51ao2EKJ1nnLzvxXcaM+WM08aJAhllA9c1
7Ol6oOacIRBhrolw5BVhpgTIHOpv47SFwvVALvGdyJR/QCwIQ1HCIOqnrLO91mSg8iecqF4CmN1V
f5k5ZmHFO/d8sGVW+OnyD8pwsXnU2on0inYG6Yv+PC+VtziNBSqgwJHIQ2iKKjJBN7u6aGs6X+oO
Piysxppb2hDsCGteYK0jwCx88u0XdImNVur5F9rPdJ9sKeDrLpgqHDzMfoBtirHh8XdshG9pOcxi
GrmfQJLHtTBSP7+1BmgAJyrx2KygAH4F1Z97zz7gxxl2N4S15yKPSvxz4mW8R7TMsP+azHwA9Djp
HKjrYijKX1H2OeMZhlSpI6tLqKoMfnBCwX2UuY2peUFwxtStHYLtmNrNfasyzpLmJwtwM2uAKEBz
IjIkGnBzny/7HgQmd0ZpXImZ9QKPm8IT6zcWLITZlOmXBvFzBI+vCpFECtikWe7PWgVQ3Mzund1N
lYKqbRXTi5VJhTxWcQ0sr7Tf6no3Y72EIZcA0P4Pj+IGFLC6cEAWH3BvEfZbigGT7RwZFJl+DTq6
gjIsWphC7IJ+MQbrgoWSV23KjA036Be5qGxyHn2dEC1+K5T4mRsB2qxr+lFa7cpNlEXc7V47ED6w
nPp83IY1o6L0rd6fphlEjI8c00Z5o/aY4lSb6SK+ZX9Wo2qlJn3ohFxotbWjEX85mayjKggettht
Lx76Skv72Xr+LjdfWx0lfPz8dXJAlYAJBp0RBkU/ssRtWyueuBOrTwS43UVLxD1SSBtd0dp/rtcD
SJuS7lnsya8NINgoZaXx4GYz/XL6CgM5pXUlrIrRKMiG5hibiRgCvQKGQwu6SbX25Y+Sb1U+tvpd
pO446yimEEf0i6OPQpFglo10e0GrCxnlt8OxHM8zqBOHHoydAFUIzoXctGuMA8P5gjSHRtcEHRjm
Y3/JR/TMoyHFshGJLCsku/nQ/KQE8veDsxVQ3fTHLbhYnEcG3cFjSV250S/0viwUHlG+BtadOmvg
HuDNc7vgdoRLx74GUbP2SmkyfjOTG3MC/Bcw7y5xveUDPK8HxsEAA6WAisq5zOWQm79k5LsT5LG9
+it0OLp5/FTJXn7qfl+aqlQCZLBzCqnURgwnItSPkgBqu0FdnuGsaiFoiuq64p72NVseyyIeW/Pg
t0xRCJF74uzS5k0MuZMAHZJvSzlFSDtJwxsi4zKDUfmhi4DUa1S7GZrZlh7w7uOo7KacirdPznFf
fmMKo6qXn27LjZnIhP87iOn0W0SVsAuT+oJR8FdxH9yDof3Jz0prOH01KytO35qth1vZ7kForad8
S1Ogri9fd3vnwe0S0J2iQYj92uGseAHmxK3bH9rSS8aIq1NDBghLU23s9pfMQ4Z+e5qEU8Zj6rTl
foQMTDo/hCUbsP0Z2Fg42GM9NwPVxAZP9xI2F8Mzc2lvLMLfBA3rwcu/3QOoMy1r6eQIyMjHA4j8
UaPqUH3GdHYPZN4GkFs/Z+A6lBxGRR8PFRxtPPuND0YOGG7pcP5Pbl46TolJyqxBvmI5l52wb1QP
YhDm4MTqlGFBfFMOuGptVMs+XZHZ24FUyzxdcvuFOyVhR6T+nxqRqXXOGiIC6AnI1Qz2uaaGeQ5e
C9XRA2XDr+jNn1cI8/DpyCmSOiLU50Zn65dEYGObZyG5Mjc/i2k+lwBQmumVqq0Dm82KmCuV1CI0
7hoOk53f+ALHb9+y8Tqsz5S0Ld9xhvD7R2oJdtF5pF0ccMHuZEHMONOEeThlDE0kz0FVXaw+yril
4qL9GtyzzQRqJ21b58hd3L5LWtr8dwpb4WJru/jH9dERff5/9MIfdy+ssq+151GYm7QkJSlgbskt
9upSjuNAFQFhIHa1QuBO0OT5VnIn81vyweCVugwf4MuYB3dSYUDP8cjwnnwrEmpFxKxLIzrzR3Ji
JcDEIP4YQ2P7lTJtWUvi2vk3Ze1Z03FAbL5PWrmIdjX4XWcIoZCQ9pDZUMzWkYD+ivJuTmGks1my
9pf12wInFcju0+2t9Y9rKNkDJtu2RVkm88tFIT6cJDlB9rcWCaj/1jWDweHC9EnRErOjrJjBo3NV
vQMQCszcqP1f417hhyt2L9mSUz+MsL06eSgqFuf4hDySi1SlzIVgWXWJVaeFm5HeEL03ZKQpNG+J
Q9iwfRHAP3e9sCr9VK3zLFKEA6KdQ++s1uOwMAxgFmplMIprfTMWeG1yJE/OEIC2ru4RkIE5/GBe
2jg1FkLgKZSSM8eiI56MW9hppWH/bJpeMrNESH6ZdVSS2Q+2E8ONAufgzDbja4DnV3CSuZmIKjaL
a7yZPzTgE6K+tJeDm7Jc+O48+aUW6HnlUtOaUA6ge+SgTTVAATKc5OKWMLZH8dH49d5S33PRNCh1
gGvPhGvJPYEGM6zeRPcdbP5oJuDU81iCD+wZsHh5cOCr+dS5aPghw80DhiOiPSYqdseWmpRIPuOD
AxUtZ/BrFJmR81H4xZ6X3Yt1zCLnUMBj4zl2PfhdPqLaXB+ZyQJ4UZsBaZLHHxzzs+02H2JhebgT
eoxm+q09uq5pY1FE+wT9JoGkkPuIME5iV8VI+rPbMFiL3sn/zrxT3vh2H05l3ZKszhnwhVbiNLbH
+fZ13PJNdbRRKQV4dVIRHfPR6D4D2TScAq4IMqj9ULHkkSbU0G66atLOYCfWksTe7WUuN76NZn97
3oA/BXOhuJQySZgd5fCoOIum1yLJRxXzqke9PxY8ryqBs5DgGr8PN5j3HpGOR/AMP2yl5JXLrq6Z
sKY4PEVnZpKBcuhhFKqAlO1rbGhRiqbYFv31l/uiJRBu0js/ASjKBjYW1mINRjzJ8XTnWFBmnTC3
uQa8Yg5fc1bZLWHHQqFZo7SCJluxEj6y8nIEnzM8z8Ezk/6iXRRZq6L1G2Irx5G09SD3xaWLLtba
6XdXmRmOa3rpOzXk8BkO8CkFpOktNsk1bdtFwN9pAnyRC5n2toUVGHXIakZ2YERXduQkWfbZ0qdz
UF9SmcVtlOVRWdo58eQAHEy6rIaLbEP5Xo5J9tF4ONlvFpBfkn4blR7RS1CoR292w9g64wXQDa+h
yGyFPKZ/9Yvv55f5m+bIVAEmk3l8hV1WP24Mup+1b4vcpLLbK7JnMqh/s5l4nUx9flYS9nYr2Fl5
uosx9yPpKEuc18TIo88QsMeIkpKF17OVC9oynJ5zN0xPsdJ50WUXH3l56y8d6xKi3zPiPjPyh6A5
CZ7RmtReO5G/EsZfUS4guMY+g98lReS91Nlk6jMohNfqUmGmt5x7pnWgO2FYWQeWQddCY6mfI6g7
2BEXoEObwqJKlO2NmXU3Y5wIFGwIuUrBHk92tF1AL2kI0b+xH+afJrhy1cdsTbxlyHuLUHxneY4u
zjlFPd4e/w49tU6+4XWNDjZyAFPZD5lL5S90EWD5tELNZQ1AFkAlD3CazN13HH/laO4dzHh8xWdb
ViZQClceLbrgEFsmonPcwcdWitKu6/gC6kJCeNV6xSeYazZ7YRbng6wA6XPyFXmAQhah1vmJSFbD
ph7nUXUEQX74lr469AcfvGoevY6ysAUpTf+vN7KiQpK73sSNXG0OVrkzDkZ5uEqS+nGElmK9dO7h
QN6hKETZzRKOde/Z5yiQH7ll9HmPXIQFhaieuFOyleIdbUFyfszFBMNrMmQdBEMWj+Ju0hMx/S6a
QTgow/490gdqTB1NFK/LJZsTm3cbdkSQPiAZqi0cW1epACVlPePmFoC3c67N8aZot5RUoWl2MpM9
3o5I9Um6dyiKcZv/17cWdsm1/o8qIEn57PTSYUjJkmxjOdDrB8iWsRlH4ejk8kirgEMWwqsgsyYF
1cpjzR1ZXaiQmRovcqSiHm6/mqWkNuwW1SttCgodoJPyoYp19ltuY5jLLZU4uem/28KaKq8qTMBl
7FjZ97trDrxiYuGYEKhbBkEnklqOsHWfT/T8kjVrq7ycWXxE1tG2ZUz8SL5HVCyr/BWH+0y3Q81D
vcmirse5EK7k0bfIMfa7EA64w0IJztBaEk026a7KdVmq+6klNjCtlg29PURtM4GtrN23Z8qf5yMo
88B85UBTu87StICf7QPB49VcRGIxF2srxYflWzHp/Zl5F36GqcaNp7UFo7qKdvygioB6jkXeutKA
0YMxgHNKyqhPUPmuncGwRDIt9MW4QxunG0CxOgYvK8Eti71VKzMmXXJBRRRE4XfDeDXasoCZbmoC
Bd3ppIceYQTCHhdYmt7d1VsbP72cIzHsTSObKUEwtm9o/kLmXQcoqFRwvIJ1gANcuGuuo7TlEtvT
VNcy8WbbzzeKmfVEdK8axfEWs/uMRqAMyBzHrEzL3GUVvlRCXg4h+wB+6tvbmM59PO3TZNyZj10+
G2QqttP2veDGMDjzFHaP4DLRS/9ojRrX7xxr1Yx1BkkTI6E6f9LH+Arig04CK9NQXcMvpXPTegjp
CoMJzu+7DzqgU8nxgZMVnoqxUGsnbsO4Yk9/HNVT67sZei0i3ag8V/NjurDpgBCq3T20DX6W7k1t
H+EZ9xoVBkh8Fl6xh9Bar0jHotNPqHmE4BZCfOOJWiwl+mhHcINiR9PBqxNIUEVntFXGvd3EZDor
XlaVtjR7NVbvDafnfWThR9XcHPcdX/oRkt2xzMnznV87HnOVTZeF4XHRuGLk71VTtuh61jmH5MPQ
rdXdgLHULxp56Fbn5NNeOdXZ+CUA+E5zpv7ZI8ehttfizeHKm5iX2oEtsdAm24Qmy/9ElAqEx7e8
s7TpIbciIbPWC4dvUQzkoeDp8cFljiEjQvWgdtOLMZ8xwb5CVcCAUX3zepPo0b24RB5r/hvcQcYB
Kcj+TrlfCBcPXuaNuy9Ln5GGuA8H+onSwqAINZY6AIom4Neuc/ns86TSJSgfsu/yqd9Jm3ic3hKR
2mrm8vuieLK0C14SmN5Po7qzoWNQ/hvCRyL28PaKozyHH+UGdrVihhY9X8RiawnovjAmycy4Cgi8
J7W9TDUNy9lRlJx85W4bSqFzlQ9o4m7fKxQhRuHmdtWWTrK7cGmI6fe+B9bjKQyz9Zjyk2NYDt2q
cgjemxizr/+CXcpUpA2FWugos09zbOzkmT6XcVGSvwDHVnD+4EVdZnlQn33xZ3bBA3F0OsA7znUz
xin3bnsxROMUkZM3DPIDzepgWprFKbh2pJA+32Jc1tk6kuGrEYD+UjIkmpJmOE1rWgBzkoPzVsXh
Rs0yVZPSmZ+p3/IxA3lAQ9tTpmKAoVTlm6BigspUwkCs9veKVVcpdIi1qerGgmnGGTUzsY+QS/5c
8vRGukLX2/h9HeA2iwwVX18caQOL9aDhsS4ZJ7po7u6xdElZVlrhEtyaSKjbCl9n6vvcMPh3UYZk
Qa19PZrzKFY5gmwXVVrK4c84jtz/g907EiIesMb7My6BtzcqnXdDVfFNUIuqtd4g8NGyubLbLJ9H
3/MgFImj95vepgmckAJAhEYmHsd4F9i6Bjka+vAMIn6KIMKqZNqGiqTXHUd+n6xpK5Cgl71OsYGq
zxqpLYP793xm1g/VvrxwEum1Q7BidG2ZuJw6LAcVyDA+28po4FjB3USn2SU4aht3Y8cPyK79BoZX
jPKK8mvskqjeAhz/EA6W2GL2rSvUBZdZVVfVRJNkrl0XHIsayKs4lhifGd+st5gaVQ2aJK8nEp5E
gYf/QYPvCYoiI8XbLDB/KThJ4ZiRSRHDN5iffW9csRROBT6uGLI/OQ+bHUgpQo2BPsJVwheWEYP+
tktRo6qgjQ8Gk/ReoOuOxF1n9DUp+3Ryx9PFJ13rAKExbBfj4iIhR0UsUNrt93TDjjEgJ1383yus
ZaXVm8Av9/7FVZh0EWVdq23fmyGow18+KFV7DC8Yyb5Tzyn/sVcDSrA1pIfvv6v2wUip2QSfRa9z
SeFK1ZEWsYLWsyKpwHCUs9DHMIhJqTllFBQd87OrdaXS/q2AnshYLrgFqsa/18My4aHqWd650011
QYTqMhZv+4FXTT40cQJBpNXT9VZJqHwZL04ahTebI4QWveJVckl4Z39Wkhqswzb27+h3C3rJfSIm
eottPu7dsR6gO2GKc+gDi4NvO8B3cP/XoszbY0Wvb8DBoePVTTIBTNM2wBqNQr0/ybqqWN1MIY5V
Is7xkVz+/tyVhgVMjEUkY442zjnh44Qt4Iny9x6BzUth2M/g+V9EcyuznmrlIdvoduSQndmkJwnh
IYLzvE1i5+L5HECTACWR8KFUWz5KfXfytypg42iKvcmARKiZKDJ6983qcMTAq6GQVua4MRGPDGeT
MhQo0KMHd/cofCzMwJXP/fq3Q2WZ29g3KZuDqGR/+8ekSNxPWWVw1zvRQw2HLRAV/7Vz9KIgYbJ6
ANv9NRJNHMu/vUzvc282CfnGvtepXEXCSEuEHRVg7F3W6cqC8are4E8AV9vHujjeAP2wooSS63JM
Cmq9r0L8F2AAHcZ9j/IxlEuTCeFN7kwnap5lTf+WrtrSX430VF74pgzEL8qogv40k2AAdaPokasA
wKaC2MslOsNNx51/TYIMBZgeGZYs6gg6rmQMrmtq9uJM+6H33YVZCTI7Tj9ymCak82Edwzg9VhJf
EJbbyVweB9Rh5kk+6VbxBKZg4eL6tNb02RsKg2RusFlPtljYgsop+kdUp7GzHK128s7n+C4RxXR5
KeoHto0J8C3VeESVrmwSmnSk92IFpsbGzB/2mx9EqFLbnJd1nbmd/n3BgqNPY2oopcqzs91gbsNq
sMk2EeqEjUnlo11wL4mQxBda7fH8AD/OPzt/Zzrw0Arj1Mxffjoqs5AzlnC7hvsYFfKotFVbpDj4
rubrUDIuQCNQSWIMd9Vyf2WzhWOHczZ9a/pMv4U7dQvwM+NkSTDitfRFdWIone/dN/UG0DZYNf1c
h6PmE62RSwgN1DvvmqeWM58vax5LapOXO26XBpXAWFUq2TLl08zX8/JaHEQAMiOHCam1zH7oLbX4
pe/j5X5mA7Oav1MmBP6FO706AXK1QJlqDl1alaExxWzKrfAqwx2wCRC8p/z39X1SHPhTk4vIkLOm
hLYP2t0ekzhMt1HbWUhoE6HKaCOV1IbBti3gqOfHI55SRQSQjkISxq0F9qCUPMJy0QJ4pAYHqLyp
WPDZSkGjnA148ph6k3mBDWTx5kgh/G2+Q5b3Ldw/OyXLsaHzfrT+RiRpyTMuo8b/v3hoXne0TAj/
CtvQDnlchF1ZohtU02BQAI+vPnA2SvhQF/y3Hm9Hv9RP+j4vPvr5I93D9vzHz3Xvasi7R6OeN5nS
Npg4P29JBFgFfyhuGeq1tK9VuRRMH6csU9pLy5NVM9nZeXO5MN/bP7Jvx0O+WI+U6Ly2KBxFQwUy
Fsmi6zjXyWl4yRxqR19FtMB7g+I2La73SVohvfyCkXIMoPIv0B4Pen8V2ts+xaYyVZ72Ux96+BQ0
XGnQrrM06Knr+pjJbQ/vE8Rbnjx4ZAchBH3PpqK28QvmV0weWdt7XdJfz7aRqub81pjy9R5XHHKj
gQ/0vno4pdyN+57F04FZh6z6ikSQQSkMtSt4dJuP/63pcZvxUsly1RBJkDWf4v9jCc67NCS69Pm+
8v2tYx4QuTdlukMtbFcEM0fMMGNt7zDR+bSZkVXbLw0tW0zgcAER9C84TwsvT+K3RrPi1EuKLrCs
B7IUMQ9DtIX6VIrx73oqMWn90Ym7q7A1THNdbBsw9cqFaDq30Z0+TueQFJTUx5GqmmxebHYDygir
8UfENpXz9V4LxzyI9Tb8n07FHAhyt0M25YrzpG2e2qci4YaBP6ElOoNG0qLXbwN6fMX54aB7G0xe
Jy9J/eNWI6k7MlBsPgjiH3FgD4/hNAcgkdooZZtXwpCgAXR66KrwYDCINQwwAH9pk3AQA8a8nrIZ
iCtsjAwE9dudj5qMMGZiBtzYaUKknuytn3tO3vtPYfyy9H4V4BP30ggA1ha9RX9h3l9x05PUBFQX
QKSn/Wm1jdHQsZGu8VnAjiUFq2leXjiSy643oPBcR12Hedra4F1dn6c75Y79DqfqYXHOmZzGtJRU
ueyoQRy6ynkHnbf2kPTLctzDJPouHefammZsoybCsk+IuNgGR9zgvIZ5ozjy2rkGyhHohOUTgqIx
iLIs63i9ty3HYMEV0nSP7UYCUJnL0CC66F8W715G/wT7duzNfTbIH0t1bcP8dSx63jEu9yVQb5Ty
v89Nl2Zi40Iyq3W5z+4a9mxfUbyeCQSVDzewKaEo6JmDGHVBgZVRWROieIFCjW/jMDXejihzOsAa
vYcUeYtmMQ0+ABUedG2KpGk2CuARyWfi29FzaCDa4egSeyeCAE/oMu+O3XyYXSCprbj2gq/Q83iM
e8kRYmARCSMIN3II/b7WG+yiMGm8uqepMIGTgSzUXiq3V9IjMn6z80dQU6HFMWsFx4yFT517pwDD
Pa9RY5PpwRStX8taCzK7olWP4cld3+7Wm3pxYSqJVCdwtLXtgZRU+wD5itkWW/8A4xIw9DDUoPYk
o+/K/RZJ8ETdyU1HF8qyv0PX/ock0ns/k3uscgpfV/Ucqscwk3R+Spvqv6sirhA+wn58wM8H72px
w0QoppvO75Lj1m43vqAL0IwUuP4gsuIvjFMrvqSM32ZbhrLSnVd8r6X10Pl9PQUl8adKwWeuR9Ee
tYpM6/dkzDqXxhQKJKbi4FKFnc2qlGxqKKBt/8IM3RshSr2YpLTvIzvvHNOiBnkX1B1/9HJL5Kuc
pLanAkhqzx5AI28dSkicmDIIuse65ntNWPnln+HtMa+LCmG614o25Cmuu0TqFhj5prWCaD5k18wO
WWH2Ez5c9D96axB0P973H0dLi6Mzbc2JWbWxcJz2k5+jybLBr1AW2XqQ6zB8KPcNuq5L+efSky8t
iQgPlK8WbuMrUss5HtahAL/rcUcGQJaeWKyGb/dMos5NEs3J8tB+xjlPVOdhptbOVEsO5eFEv9cl
SCyotdy3F2/wgzbHwgyoRvyjmIYLzF8V1yXw5kgAx65/18T8JRVcM6lWZ4BCX31Whn9ZGArj7GuS
208gxv4aONZOnmVWjMvRPhTM3mlvFFy5UKQTlFrEFLRmfw4OSal2FHqKYL5Vx2ofNcvtwZcx/bRz
FL7UkeLKPAZb8Xsf8L0rAtbJtV25IxxJQyZG3WOkQusw7pGYq08+1f+bFwn2UlbFVNr+QAkwwR9N
boRjWGfG0os9E56rq/MLH21D0fFQbIGZeFwgtEW/DauqerVyLnsJWRwvF+Y2MWWfL++zfDOQ9QTp
BpSzM1isUOhM5RZ267M9yhlhtGcCs3lrc2LrsOhxMblA5whmysTt3HJ83nIv9rkN2RIiFWrQwOis
MPyzHJpm/+dL50jnYxpxxBgvq+QabINFsIrR+qAX0N2hwOGeX59C1eQxwMgsYnYI3OhSPlvgVJT5
xyL6CR6+9Q/OcncB+bSLyKMD1e8Obbakfd7itc2cFAyBkYIWvwtKPKIj92l2FiDnvE3KqxhzebV1
F50khxxxZYIxGcsHWORvoNzs6ispgeb/n/KjE5fk1NzB4w6+wvf6/VaDf5DI98WVVgEW/XwhRIEF
IalSbhaz5MTAO41xQTSAk7t2wdcl2wsn8uDuDYJ5n6unqpgD3IBH+n9JP7JUEqAoyzHb0oBxEvGN
TlYczwwjxtfmZpjp76XoZh1XA8ylFDgAFnjaEgfodJXgUe1bpiLIm8Cvo5dIWTlZmlPUge+a8CRw
azmIF//yDITo6Sr5wNbuVUjlEhM+nZUFYpS+7W0rvJFC085QnGdgfI7XnUGuUQbVlz5NM5Q3oCl/
ZwhHB24jDVpYqMfYz83cVgydsAn+lH+xPF24Ko/Vx0AMyacIlHe53wP0eiSnmB2ycqf78h2BE7kQ
kQUXIpjnHuCuSpjBvOPX1vbpbwPnARBlFPOo36ESMLZ9SqAvORgtX+0tybQ4CdDZWbvyZDqooQDY
PnUcvAd16/9ZTBS7yY3DQHkPl+0PJPwclAE4hFrCeaqi5Q66p2/F6vuB9b1musbGU720ErBsf9vw
kL9yUF39HNtX4mSmlfM4nulHhbwJ222u97ta8D2x67LmjKoh+z4ilwp9jwm2raON5qVOrIr04Ip0
vGP499Sl9fE/1fBS+YOlm8qbEgCX9FcByRwXptR2QuBwHLyewgBzKJPW4AGT85kDuse3LNFDox41
bqFxZnL/v+SW4lfQ2nw3FOapiQIympzGDQA6aab+OdEcLqc25QNShtWOL9IWSZygok+wuWw7Gdlj
S/IL1oewrt0lingW9tEE3oPRYNJvJNMg2dhXgb4u+xcK0hfUQaTH50V8cjruIeIVQfLTDvdYaknf
TDLpu3udk0dr6S5pOZuMhgUtVfB1xkczLms9YQK9r77o1S3aorTyfLwdVZaSrn1kKt3MNmnnyZTx
krQ8c9ChiaN6byCcoCNPCt1/0qGzL4DjUrErVOAgjVjoVe7tK8bJkGy9m5XAmFKkRsFFoLoh9E2q
AbnNg8E2BcM6EpIomUYupk4CG2U4QkRM5FMwr/v4xna7QYzpTK3jwy34pIXwrBx/DPiAByGjxyjC
Nc2/XsgXQj5G4VjzXnLhfCu8HbsrSpw2RNLas+ouwLOwml59xpVdV77vU4TQviwBRfzvNw50HENG
nxssGVhTsWb4ErQzOg5SuDbY0B99UII/nAjOhV7n1fcX4Bso7xlxD/a4kC7MKa19kU3kMviiF6nr
FDnxktCKTfzNUYLMbccP38OPPEQ0sC2RWzFNQUlMvO9Nd2Q0S2YRXxL04xG65whn61qYLCBC9Qno
VPWHEb4QrOrupKfiyOrNeaTBkoGfadMhq+AwEmrz6Crr/e9ybo3cK7Pftz0gTK856sfroKsraich
y5oN+xzO35FfZIN6O8/q7Zw/ON6wByufFsWM0Sh1hhqHROZP7s4q/zz3nqc5WTsYYlZK3UlCWChM
vFJGA64djpvEdzGRz4WNI31b0uMaiwXzj8HU07vfd26qRLn0h0A/WRoEB+qcLXno+N6ENSeu+jbT
tAad77BhZBnjg2Nwj5lQnfwoTLsBgVsDlv12u9PYkHwUEz752R+CN3WQczP+ovMJ7oYGGJK6XFAP
QkmAtey01ef8y5hhtEP/R5fzezGDNmxa8HmiDOxHYiJphYUiXz+DUMaW9Swc1vr9/elC5iChpamX
p+GG8hRERrHzHrHpdol9ZQwlzXlacodxvn22vjKy8J/0fHbkdcjALF5qElhoN4B7cAbaRlo5Isod
sOklK8esu7Pa1Fxyr5GMnDOacrT+CoMVNnoWMlTxKJ+S6fMHy1b1iwjZcEsz7zlrWOb/9gMigDd7
WGniYSM3w6c2WDB6tO8S5KpFVBaORMYj7MEBvCKhvENctHIH19pgk6kVluJf1TNDZ8SFQzAoCQKe
4/V0XlQ597td0Scz+F3gaZqF0Zc2VS+4aMg/xka9FilwTDlzyocJ8BMsyghCBhr/oBVosFgk63LV
k+JnwhtVkoNPNWhn/4JiqCWJ9kWapE//Dqg6+/61+9AQNe1X3W14Zvav2j6mv1ZgyIa8eOR66Pho
4lWovU2uYSIJgwLhcFGldzLtlbr2Yy6eQiDXwrUTk/mIcPO0mSP+3g79BDc68YWzKQiDCiTO3xY3
kMR4/enYlE45XDCHPvsAi74vd1DnTEiCUj3IvVW6/w4neYpnr4f8sOgMZDkwtdrcgfzq8aK/GH/e
GJ4oBxpiQrJk4OR8j1lbtVVOL4YqZnztGtN6m4Z8iun7G622nJD5znUxLVEH05cS6dhyZKZEhyUH
0oDwG599338UlRkltQCzDVPaoImZ6IKaMBLVFaTBYeFncherzICBGA5lsL9FlMo2up5iCIKO0tv1
l+y5+BD6nbNfsdeKFOtMJKaYyuzG25w5saMRwrACu8qjF+UzBTXty44BhYWuEBBIvxEkd24Jw9nY
4+jdbMxblM78MxKexSGFDuqpj+iTWAO/EjLWN3XBU7dSq4WKP17AY4jKkhHU3jwYRKj99+qKc3h/
Et6usu31Ull1Zv1rPzXrZOr4vVn+1IlizBdr4Toi5yRcmdeSv3xj/twSR5evrvVmx75rTCKP2QHi
BGJxkBqQMntvn0EmDMkC4h7klsyBe3AaR9Wz9wr5akTHseYW/uH7BAvOQJxJX55rPzmh4WzbY12K
4rcx9CUID4gug6pZ7wAu4eX/MCwNwYumUGvy0geLbhSFZAHHLCsq0dFj42jxMV74s8CgCxAG1X/8
iyn+QK66dLIi9VHFfiCKYrG9J/k49cM9B5G0hqFxUoQ8bcbBb0zPbN4Lbs9rP4saHckodxgHvi2h
avqd7f1Us48lJt7MX+YzKmv0vhC9VsoPQSIolinJiw1tDwoTF/DhHpT22axixpXmAv9IMSXhdeI2
ePq14PZdmx/KR8PripgIbEtjuJPDy9FuaWojEZkO8m/sgYFAZR6mEB8qVlbT375/ECXMdfZOmlJh
n6abFxl7zxHnmecG35XiwC8xgaIDj5sJEQZhs/jbQ0VsMs05K+E2iX2e0d98UzOe6LJNSmW6ZFxa
Nekm6gnxoPN5LaNHCiz9rOt+x+AjUmxkst09XXFjzs846wRBulxWSSt/ENLczVFDDgDCRaY/Ba7h
SRN3TNsdnIJzgnLWnNOlECl81QBHx4n3G2hPX9+mpkdtajWH/nZZ/ulhaF+ld0gnKsLqzUAh2Pqj
5uHvngyXwu29cLAdZAqY7i0SkJ/zue/5bB+mZS0RjQLvd3DrM717/e4zSmHzrELpajsARbU9/Lzr
3/tTQVHYecrVM0RnBnSD9cRFis2yTz4xC8lgUq4bvArp/dbBXW3f/KIgT87aywjpltBGCQuACRz1
celCzdnlsQQOPRnOtowdfy+b5RJ/OBfcbfafz8JN7kYJvrCEx1pzJ3Qp8Ulnrl3DzC2qK/MYdjs7
r5lMxFh0QRZlSQdkPhuz9QtkHgj/a46gJNCdWej5A99YAe+EOrDJS/mC+IHiHpfTL/xj3UvB6LB5
U0Ze9syw63yRXfhkyk39Gip8CwYffH7d1307dfhjVFcGufyO210pF8zXXrFPcNVX/XAkecVT8qj2
omFFBrAqn1/LgODj7vrMZiZBj//sDkBw+e63+usxCUL8Vua+oCw02ApT/kCYWSsJjJQNU8EaX0HX
9UGC4imPUCit++1ovGsoffcvBU26BlKkJ2K6a5FgVyEOku10OGQzz7BBcx2Xif3ICx0gSx1U/42V
aakDA7LyloZCWNUc85gZtzUFVyB1EIJM8swXKDKlgwtPa0FT+5kzWsEf/D1QM1q+6a4VY46F/T+d
XNNwDe6w+WDiT5VkYcJdiySC3239QOI35Thvfp2xrBFn4PohEafa14LjittEHFEPNKxhc8j9PU1h
ljQ3Cyqh87/l6upxJoUrGUJpv+So0/IMMsSThnNYvwGawYhcGoOKwcyzmAEzNPXEBnyoOrFRUTiR
3LLMb3ix6ZmponCw1WkE7gPRTipBVlpZUGW9jzYgMs4xm70Hxo329XgeQlkxnVLYKgZxJQP4mr+V
Ed8bId4geA9eOgosI4BCBXaVkLFmo9E+Yii4mJQMy2xHHxYMwh4Uo77yru/9L6XJ1lvr6/d3Wfv/
GIYUznsnVhL6KZpY8AxZ1QiSY3PV5qvGSARift0IkyNEp4JBhf05oQAEwOlher2ALEsRqZylEcem
VUJZ/9ENap2KgGidk0Qqwzc998E5H5O4Mp1kN2Df6HyRF3o3UQnbMq2VHcF1UZDetA0/WekEK3Kt
51ETt2Ijft59Tc00oTirYFXv7Ac/w0dLRBkANaIqq4/BChMMXRunmir/YIf+ujVmLnQPVE9Cy/K0
nIvDD0eLbMobsJjMgMUFea8QZaz8qOUCRoauJ44hi5qFgGL0N9cu0vqFmdQhVnFIAXn8XoARwaGe
Al4OIO01ZKk1k08eArbnOfpFw01UGWVVYJqML5egaSvEzNwZwD5/AVyIdgBFaV7v4N4Ui8vYp8fO
KFpbD8566F9zA8hadZP+2+AE/1bBzAx6wFhZcqs+Dnkv1c82h73XfeKhwbhdRMvIaaMJw+zUNOmo
9L3CrQ+YF6ptau/d0mhQALp6ZN+/m9wed50zmudOZkVslHGBrfqlC7Pm0Rx+7JRdKG8ySN1C1Tau
ov8ZymD13qiwVmPF5GXMEMhmVy0Dk/Ql90kKDdlKoCAC1XY1CAyaSLZvG0TWV2kU0RVNFCImmU/l
TYyH4dyxtBOyytQ+tPxIWclc+1F32UXP/k5AuiBvB1wOiTxLlK41lp3jBUi8sy9l54Qb5CeKrOxV
H/EWlg85KhptZODn7t+SeeWtBdSt/AciCsKWuFUlhuq+E34SGWX+W6kdp4UKr22vz4xdYUDMtySO
NtmAVGjuyGtYliTuVt/lYA7SD9y2BqWLD1Tp1Qa/qORvrCOm8FYife3IW1q8oG8RxKUMEyfk/BCg
kC4ACXSYfPTBVICHWNUapH1rDXQeRYaGDdNaltVi13zbVvljAyZ3BQgMb60l1E++Vurk9JHRFqQi
dfu1T0sbGB78cMn8FlmCnbQRgrFGAUUgTKWv7TzIA2RAQQCnYCTP5Fh4S53k1/KJ77jvwQmOk0zo
+U4T7lIXdfGwJm/1TEPYH4KSzwRsuEaGhaeiRYMcqIx9AOJNljk/8uTAF0EFtmOrliU5g+CGNrJc
GOHwVBzdWZ0XxjG0P3CdBhQoEUNKtVXO0C3LvfFJ9zLbN3+DaGnF1iV/a2xvN81L/kGuxyJRCKFb
aWLonLeb3ZwFhMYvg/ROmx3qBAH74eG/kOnrNA9Yc1kLoUCxfZiH4IoAMPgIvWryzVUL2WaiikvU
lfEMEI/3dOH2HWE5J1EFhfZ5dt2y53fNkRO+r8OdYpdXBUZfG4rGpNA6l7NzSgbmwpxSffT4dAvL
j2vQU8K44AacdembKtdAmsgQ1ALYtreWafOVurCn0PeeixqqYhxG6xm8PZ1kZrnWwrlvgKXTAXMz
NJg+cCDIymlTr5JZtrVcAmo/4IaoUiR4UHN0KGwHEm5kxy7VhOcud2cYsxv55G6pGc2nlIYbG7Tb
+4GHpdssaO1iC4AqDyK/M+acJxRcM/B+JOE/vufaddf+aNc/sdGrglDDNawg5ir/66eHi5Zn+mU5
7m3Kui9/biPQ3r8YV3QqBTfoHR9qPJhnF9zP7dZrX6O0Xf9LLe+Q7oqxAFEssTF6ZD53VxalFF8M
qeO8ONUG42Fjg7gn/obQzQbMO5LWb0tWLbRcUyJqvy4PeKMB2Nbeiwf/1PBcufZHaxGZXKoRLbmS
WIb9WJgD+NR7chyXh1snFLQjaHo4NTgQND/l+SfS/F0a98Whj3TW4AwW1sKsKZ5a78KMfn1Y3Eed
GEbp46n9OYDyOPDc8v9vUrYPHKJuyIIkpo3VTWrqFq3Rp3GDpZQsPTw6gDr61Us32XpgFmm7MpYP
BucBm4hkV6gGqo2UEtzbHCioBaRuQyRcHuUZX2OMEDYVF0VBX3kBHm8GpPdw6EBARbe+fDn6+4H8
EJafCngRr1yjf3ZOw6xXeDtS/UOIQUUWtCv0aWM/pN2GSkwWZmtYI9eK0vwxSVr3iGBuzqT4y3J7
ZU80hgZtPwErYh7wML5a7KgMBHmOoUMJhHFX7k6ZAwohJXOGCmQTzvb4FZPZc5NoSkUn3+Peo6Da
oO+KS7lOsXremu+L6fG9TLA02ne1+ibIBM8QentIM83vqme8F7NfKpf5gLs2aOGSe+kyT5KMVsdA
S/WTtzacZPq5lMqqL0bBN0QK6gNh9IuotMq13gGAkmzq62dc5/085uUa8hsf/n35Kdn0Dg+6V8N4
w21T5oTpbMQtLsRx4O81e3avwjddaM1y24iOwX2hIRxPW24Qq5/PVuxvjs3smyOrTwhMN8Fm5uPk
nQZ3CvC9Q3K8UeCc6LGRsJQ68XeZ0t4mHrdPSASaLZBFuZP4dO+DgluISL7p8iSi34C7untPB2E8
pgI5879DPqz/wZ9LH9m5byG/jH6vXPhqBlWHddx9PlbEWA+owLQRZ9Llog9B2bZOmIqsA6zGLANB
NZ8OaYWVUbklabMXw2eHqTD+abVwvgVc0ulcT6TZ+Bz6YSTUK+SH2xbK4v+dzyimEbQy2quG4cjf
3aDxta40nXy6qJawFyecV3HxevaOspnPB8m+ukvB26iFMnEqDvVlj0FLyR5zVf8ZMfHuhp1lcPcY
EgANgrsX4QxP+p7XFy0vuNL0uvhx0IziuXBcr/S1Niha1iFXVmplHORYPyQGyXQ29qb/FpQZ/Sbh
glPGE5oI3P2LfT0KPiADQCfyJ3MEI5bioNOxcBAgcwg0CMN0OqpELNGLLmV24AGTB5AkRBn3IJmz
zcP3/JmoQ7w6MDNPSEECkeGaKLbxzHa0r53aUBxrn9wSTKbKU5M8K1upX5oKd8ZmjJBnTvMul79Y
zhJdqDcIYqSlZe8Psjxxj/+1p7v2KbQ0kCh9L2QF1DzP6OEwpAMiT5dSU+Vcj/tD3llYLWvzxZ5V
APzxElvB1wIToMsTabvVUz7ua5LI9e25MgTlX1mxC/rgEOB2L1FNsAHtWxa25CeVyUPSXKHFu8Ab
TutPbC14clWv8p9qG0/CtvLDwhzmXWvbmNUfp4qGosulUMMP2XjBhQDkjIL8wd8VH2jDvR87+mpJ
pHJOrG0gXGPQD5idYGQ0TUkd+f/8DaXpEFaSijgMsJBq2a8kyWUQ8bQWkFWVjnbjUyfRHFF2ilC2
MYm/VTbStbxiZMOs5h0PegfLN7DjvUfaGqmf5TlUOT6pPoiN7rqSEjbNcrvZrZJHJkTVh9A1iFHC
bu+kozMxLneHl83fWprwjaoqoEy581amox5+n96HOYZNaIUBYWbQycR0Zj0rwtZQida0/LAl8gQu
hf3Gjh/Ex2zehyFLpeWbNahLcKfYMBDh9cyEqROYqNysvrwD3vgdBTDbU69GaiHrGCTv2hO7UDxO
CTGYQzaPvlCMH1Lxq881iNtlK0SgM1YKjxZnqgumpa1322hsN1vlhMkybg+52hvKBILqt+5eBIWY
pRy1lexkEVS4tCc2QrlvuLE5pTudIVCr6s27sv7HPnJLPK6pZ732PvHZP7BLHXagceM2yFF4UDw+
l6qOLn5GoT0kIHsHI1zZV9aMP4SpdFl1OSApRrce15JnLDnxwh8lDwHTXi/ZjCtbso9OGipGWHWB
qZKOyf0o6fIhd0Q8cQgSs/m3ezMClZYc8gKJGnU38FIRhm5oHSqDi/htCa1O4e3QS5TZyb+OOU0I
/Bgs+xLolxOFI/JFYwHMr9c0/ssJ3KLDctkgOKApWgxYNQGQIEd9d6VBwzwjr/qU3CFiZSuWg6CE
oBzqHyMdO234xK2Pas8+VhsnjffH48ooF/wGlZC5Bhi9t7r7YC4ASOxaUpkh7Bjf2EDdmZbBhDot
UVu9tLXlHFV7s1Yd/m1raLTR/X8UJP2nfVk/8+Ux7Iq6ZVdlj7vkjEPkJw2dwTWOx2Ftcf9R62v7
3r6z+U8sP+qccif+3fdWuxqL7azzeMNSJvv1iTrRFje0TGw/guX8KmV10lH23NO7R0Zj1MGfHxfS
KUjV/AYeIJEprj2fqMGmeYQNEFInNQUQFaHSqoYUdOmJRxt1v9zOFMEhz0AapsrEX5AEWTkmY9qW
AlL3ZDj5amG97FJMwta+q9fZ0knkfvstHWgmPzHDQYSCAJbbgKwctHy6YSccHGT9mme+Q/FJz/+j
iolJ25aWBc62Keb0pCLX3JqS5F2WmQmnEoyEbqheEUek3lC4xTxXLA2Ni8m8xkd4Cq1o/Gr/6XgC
9IanK/VGDK0D0lCTD9LVBuaOO73BLpNcmyfOjyaST3xNRGdHrn0wErjRphsGBZ9Hd1hvnpVndolJ
uMgKbCqxVaje0e0OsrjZe+vl27oTr1JP2FtW6IgiTw2GZFk4q2ZYosDO4Wwx/96CF6yiwkI3MLuA
2D7Xyn/asqqeMD7TTj85gH6r9Yuy5uIk/VUCG/FEBrAuxMeVMCqQ7RuFqGCfzs3ZyZOgbPIoiD0n
7TFa6CTyNodyYCgCfcnnI3XHp7NzhyauosTsTUl1XgFpewIZe4oI3d4OOwc3mxCM1gVpNeovb+Qv
v95/hQ6xLzBnB5sFfDtND2Y1Ji8rE4GTYq2jU+IhY2VpBEyp9wZXEWkWDfon47ZVqid6UYf3dx0N
j9YMBucXIsRBOnklqEXBGfOIYwCLWrKbxQNGQkMPqG8izBif52KMD4p6JqmhZm9uGz9HStU8maJv
2s727wFRphWpKzj34bNF8bft2KE20VgkmqWTwsO8GXJFzlejwmGBlGIFybyx9nzsKd36pv/wMnwP
+qkW7eV3UxAefZe1ZBIokKzZFbjJiXop5CuIZP37/3smMQHqGePsKizyQJSyCG5VM0FdkJ/k1kOm
LAaYeomJR+/F9OmGB29DUGV92SQvaiD4+08RrxP/oqLhcU5+33eBbG0ZRgyDictPntsCAeh0zQX8
1phDBqo+RUqsAHDzoGqlaR6b4ahmffk4W6PlKcJpmrT9p7VyZpyMG1dRmHj6etZgZlxfZPnWYvmN
I7TyvkucQy4aeGqVudEagI4zPKk6F8tkxZJRCPjsVsSe2k8anLZqWyG7fFdDCJRHxuntUFXnkDee
XJAFuz7rxw4RVaFQoHvZynT+b7VBz78fE/0Vtb8b6H22uO0ZOA4/5qzRfjPrh/dSFgq1tYbgmso/
akqH0/pK89HlBYtZgl0pvIDVZ7jNiWaGVgOniBxejIYUWvRoPY0HyS/S8YemiuZ40Dw5DRvZhKYn
3t95BtpFRMahtO4TDowEi9nOCu+HKhAamtmv9GfjpK7eJQ/TaZAOnN1/O+9pi073XPuoThJSuQlF
FNpQ3q3/rpZtV0qyMvzHr08ZyNPe34MEsUkqLV5P3OCRLtSz930XIO5e3NyxIdiHRx1gRQhHAgsL
KtIDmKx4uGl6jbiY8MXl9MkTWfytM6TWHt9f8wQjiMl3rYhXYiTLPWHwDIBkPLuh75JA7PMBnwtm
rRIcobRrZd/p+cfjv5CTvMIkRp7LiQcIx8Tzg8AOZ+W2y9mpyQ6uUfyuN1cIpnBdxSWZtVEPIDtk
Hg0sSLsUHgVMJpcJCwBltK+sUI055f/QhrC7Az0z+ATlOt9p1OcRXxKag7tMZHiGIC7J7sbBS598
dvmCW5fNRehXdhRvry4eO9eLwsu817Xy2TdcK6cYSGBVe3ZS0FgwxHFoaLkKvJ3NrAPwAptWBrOs
7DwTvDPuOkWJWaPktvkNYD+ngGpqmqYJvvHvRRC39cAH4OjPwROle0BLjw0miJNjmsakpI3YMfo9
kCJI3ZvD7I+mV0JI2M8kzuzfEY8q3yhPrXmzPuUWJliLmZsQqZm7R8f9u4QRHBFyqip/VEPm0gQ/
7jGOyTsuxXi8I8JsXfI7qis66e55qdwUhU/Akoq7wvZrfrv3eJyxpMQEeE2QNwNGTL2g5h9WvwAX
6mP5TJRaIJiB//YVi+cu+jjqzQhN6D94r1FD2H7NZyGAo3E3S6Bw8PCAo/nAm9uxiwxrC0DdUy8f
jeKFaOku35F15QdFo7mFzRO5Dfj/nodbANhkacQOTnDeBddPKjDxnuWmK0LAhFRUWb037WdXFBXe
1Aat/C3LymQPWhv4YBytOSqhReGkUbgeIW8XfYU5KfYu9bBrF3bApuk+YGvxxce3CbSmwRXS0LOk
SeIeAr8X07tiFg/rxAsnp7qlTqnFfbaswmDz0kAvrCmCYBTRun6xs5RatT/6boMEg//5VaZ2G8+g
sa8P8Sn+MF4rgjA69rb5zzoCdBJidf6mHvpORrQ8w/9b21Nt68p6EIOZtKdVSiAMS5Srg1jQrEtn
rou8kCqRAxyZgN4z3giBjH0+vMJxv0/oWm4IYc9cOOXEAkCH35S7EfOASQjwy8yo07WGxKRypBm8
fFsB0DCN3wz+uTR7YG6MxUti8RtJD6v0+ou54Wb/bDlzjHEkXjvprPNxMRSQTGGxYxuu2ysmH6Ve
aQW1AVaAp8XtQNhRQU2glGxlT8B5liGVCC69o9DyCqu2xq311+ey7J1PCmJRnKp0Kgh5m4BFyedc
PBzNqWOOAyy4y5hLn11+b9I9G9XnoH8BNJOTj7MrYP589WYJDluQbhVpflO8WpFL0FnaiJeVERBh
GH/tKi7NMn+eMu2STFo0wB6j6+aiRfEseNuRR+GkQ8RLnuHmOvyfGuAlCLKKzuxdNfoRuyhcCWny
NHCuifx3MW5PxH+ZhF3ZZFb/2WNrcdvC8eV1SjgwSVGur0/WI/pJkHtnlS/zAtWRNtpWyfE22Unv
qE23ayWjUoncaaxhXAr5tc1wS2FQeSONMSZUZVupg1rJ1oD+Zvk/BbwUNOPVv4Qwiz3UocBnEtba
r2WNu8vs4IBbHv2jysYchjHJxRIe6PuQyAkmjzE31Fou2Hjr+UI3gbpysmjicJwBjpdvnAdOE/dJ
kpHqSJtdSkoFZKndtr0MSGePTeltsOoPCS/3kC0rmYf0xXj8pRs6z+vcaaV+7kW9FSQrgmAtKYwb
8bmXZWRU0fHDKEMDozfO4VQGuZH1nF7fy5p8y36/4QvYqxzma+TlIULyPcpJQazE0nNYdTW/IPXP
9PKcBJX75cfDBKDhh9H92b6qGRdTmEowxU9aUStjq8fgc1r+iSD7QhC08xZD7LdretcNG0OkIogl
wPZ+t42PUa8fiJNJ8oXg9Q9a4r/GUGIkByilwGlU2bv4WjYES6yG81TYNz1nkQOmJWV1sA8fxy8P
DGz1lXM2Q0skpbfo2w7U3VhDxzsEmdB4vP9dtgwg5Tp87VTepPCN8hoJYrApbPeg4gu12yi6eEZn
zhqyHSkUv1xHBqZUUPVNDk5GNSCzhnqav5vLHKMoZFETw0NS4pP6o8sUVPRbiT1YccapfJ7nJ1OT
06bWyQoJIbOBDxGWxvqGk2eYMZ4RfhWEx9uB/Ia2pMhM1mzGf4cBKQ1/GGy2sKFUmZeSUBfy20eo
ubbspcaZtIZoasC6l0ulXKHlO8kB0VP21EL0jJgsW/kIge8FWQo+vCBB17sZh8GNSTmJ+76QzriB
DWOhEZnYJUvnXJ7LVze+C6+ns6bZHk4WlCbhVsp5XirXoGKjuW9nNMjCk5nxPXcxFW3HyOawlfeD
/wSiwQKzCwjhagycsB6Cy9mR4aIu4/vL1qYZeuplg7q7Gh2xHC2rIGWfZVk6zFZTSbJpPGSC3hSd
Uvw3jM9puUReSz4ilUwey+fCCE1SgifeNjjPYRvZM4PDZkI6cs2oScoEecvWgbZL7D057wjgNjQz
fkMNPxxI1dQo+ib9pX0u6Su66lJksW5cWcocEVdGN7n/fJjZPc5OwhrG0PvkiiJVrVLF9z61GmjZ
H4VIyntmvbcnrUBbTb7BTnZlxBBKNcOAVfXE9FX6KMD9RP0In6S69YA/Yt+QdnlS3Zm65wlB7goZ
y1cXLzez65BK1WRaowCCRUAAOPTH9Yo9n4jCpJfAc7mWkbEPXGQSTNz81WwJ4rFfkubehIsNcm3P
nHXDfTb25K0vuY1C52rKO7hlOWmRDlvB7/UjYzODQ6KOf5ErsGIHA9CTeLI1jMMuD+UqvxVYH9l0
Pg1fUf4l0D/k5/vQ9UeRrVWeg9+A85nJlgK96rcYO0QHfMtFWWc4QPo9jnG0KnJu4f/WZIcvbXeX
zCo9k0rmgjl3a59qVRMv0ZENd60WWhChfeaUFqoajSlm4PVHT9xXK7rDk7eIgPSfBi/38GiggBLp
5SPMZCmB+I7H7fwF1SCnN8/dJw3AGjaeusScNMiI4gJXHwPQgB5yKkAAS3qzUYmS4mAoae/9uAAq
OSVukyH5w593otUkrIGjzvrMMaIgHdjJSRTJbEF5ZH+coR/pyo9ad4CxZPPwMAUbkSmOtZiF5j1O
awEtr3Tg0ygoPeA0KmYOWj/M5Og51LcFba4d9z0WfrpQ9nW/Nd04cZqoMJjnrgTV328Aqv3EoCJO
phm//ZJmvUm1Fo1pWpxHQz/P8xebmDVgXXR9eQ7VSn7Rguy6+fJEUyF+UhKobZVAyzURAfiTou7M
40fDAgAaStlhRFE3ce2jSWP/GGYsomLQhDYjN/rZrpw1HpfA0ZLU2wya8BKCgETTbD4bGXgetRvk
Qz+w7ThBm9W0D34idFM+lZcHvI8qpwgATO68d2y/HC4z/EgT7+uyWLI2uAlq/YphcwVv/+NnWksc
gRXznOWueMU9HsP80vysfGcoDH1WcgvDfApqrJs9HcQZMrmwn/nu7a1OFrgavcjusFNM7RyVkun7
I6up+U0wWJQaz2dzqoniIj0N9YODuBGUOjGXPHBJivm5uGLVuGWDGHkS3/lYuGbTUafif/QqqPT2
y72J3+safNGWemQfkKWEoWjusjhLl2ajzuLpDDjclZ7jd+IJugk+CAue1WjMfCIVojwk/b4VbjTD
K8gZOW3xSTlBUr9FdE9mN/VodbhXcjIje3pMdla+A+wy8dZiNM768yeMfJpBbxZqbOteyox8VkKV
/QpnLNeoIc7vguBFppZasjs34HBabHJW5nCIUuu3wV7/+6RmqL8/tzIb3X1QXKXTqgMRjaQAebAi
2wTAToxgjmoQyq6kuHdDXznIiP9XPCWLiAvBs81K1AKw9DGpF6PlaZZ66JFnw8AqHUaykVR+7KP9
ie/B/Dtxx35z9Jf/vQGHVshsb6JQ/lZm0DutD18exlQAr+VL8F/U8aWa/ncH9tugYyEp57tacQ6V
Z8VLSRx6RKcrK6FvY1gwQEvH6N8CV+X8fncz5jK9tn2HcUz9FKngmML6CnquS9eUTAZZazfbsg/n
pbEahoX5UPk0j2TyMdAskUSDc/sJW+LazRZvXdtPVPQuSXBrxZu6U4LTD+bb7nBroqNfQG6tqb1w
KR57x6ltOOfU1XFIUiR03cKhLyBC3wGq+kBSLo/xmjuPD6gJUm89QhdmnWtC72HV21VcTy9r1eUh
a4/cN8UpxQ0wFu2kIeq6FJrHEGyNlQGCA5+C2ozGFvY44x8tnPCcgU74+H4aH+S7qcqg60eaUYJz
1dZgPvnAJxC8VE2EeVSsnDgQKcV/F6bqh6j4HONBykMci69exxvdomqE4JggLYF9x0mtFWlUxd4K
QO6RspDXYtfW5GOrjXMNeIILyJyS/pGINMQAvt/ZQ0v57taBGviHcd7EDsjrZ/rYaeuVy4KaRp/h
bS/1xdbeIcktYTT5ai/eq6h1rweR7EommrITMHnexTlRAf5k9AnL5AD+ZOlRXOfUFhulbeRembIg
AUa9f8qPo7b6ezCgCZA03w2m85NdKL2Munln0MjfAOr8ysqxnWLXJT2XDJfCAifWB3cmPEFiNMGr
fywV5DIXp/4kgST1lQaPDy2ulyEbE62JfPlrvkycJmWj+qtvnh4yzygUX6MihHmBa/E68w3I/QUa
IhDUrPT68jIhR3UIIqYAxE8OjkzFPrRs3yobWtZWNEMj28/vl/74F2l9z6ez/EdwZv8VPq1DMBbf
KB7N0TzuSpYo94YT2fa2/LY9VdflBVaJz1W0Hc1H/jNK9aL2zTSdv7izmKSiReHP58FP8mXpTjEw
oiB5bytdfW+NZ3bU0UIjJsjek64czcPr97g+xekVM5DEq1c5lqz8d99cu9HAW3B0dHcHeLJ4JfqZ
2QHo3yGDY4enjKoVuJfGSpbYz/m9712YHS8HtWbDev67L7+28oRFdTKj2Z2Ox7W16av+IoQbryzU
Y6taOzMgR2maNd8wFyR60FJPxtvxCfU7kcxdbmzQFhhUEEUjwb+Wsh0KUpaPppGfqpNaQSALO7Dd
YlLdVcDVxpfLTITKb+cUFph3X8NtSSvuwrAK1k+XrxwhwtdEEzsrnZNYRI1fJ9EsnKhQB98FOjW3
Od0bX3osaM0Tauwue3EBSBaoXIdXlwuLYGimT29mkXhcS/H0dx7yd33KDrErFuSGEptXMGmr6U2J
56YSase2LYEwzQV9tKh3csvP4dYwLeKv3mJZMycxBdThK9ts83q/xm1pz0bLpOQNnXQimCmID06Q
YNOWksvsXg+DhNE/f+3M1qQaLUXqQG68dfn43pCS0JgWjAO4lDWOlM9bge7vzbAj+K7iQUXDPk0w
n6SfIcL0ZvlmQL8l5Ph1PM5Fl0URDVssV0lsCEQBqDQX+YunwTeYYHG59ZCQvRGLGNj6kB1zMzFX
QZfliPW6NuhNKMINzf3kx+40hjhSlwxa11vVt/vDnHwI2ag4wBd++vfYXTeOzrnWEue0eUN2xXZ9
Bz7aUfVPCotAAMbzAfHWjIpLfjJz+6TYQIaT7hdA8l6pdt3eBCg7Y0BY/iEAY6nd2OxoWXBIwZzO
dYJYHjfRtrigfJ1qBvaAuAYobHMeaYNP2lGUsZgNGvZRjSlzF1c53J7u68h+R4R6E1oYylJYzNbj
i9T1ClHWBibUwc4lAL/qX4jiRCcaVYQv8Ml1MK8QXwXP1Y95HUxYqfmtSGIawR6tpVTt+9+36eGv
hjgMOhY1tGObbuXrg0rzCAxvl/mUm5230JC77LagNsPO348voHyjcxjGBnJBd2JBZWnoX6CGF5Zt
48m8STitBYW/Mp1eim6ydRaylZSSw1jD3+Upqnc6ik1iIOI58AldrDlW1cJXiaXiFSCINPpSP3pI
CD4BM6cgT/D5sZCQ+iNtOF902hJoyxh7OJ+T0BBrnaVUUPqQ1GLNyAJ1U6WSQdITI1WIWQnLXjwh
Zgkd2H7Gb1CByd5d4aJbBVTFgFKbb1xIH7uO1ORNWiy5aK977mv8JynqFjWbui4kpVTrMilTg2Iu
jMay0eTMMLVGE+EybYSRLJkf3tmXanCEHx2d0Qp8EeOc45q2rPnz76IAgmMiZ3bRM6GzB+k9vUU6
F8BiGk37D6SELcc075WLajJXUx0R0zAJdqQqWb5r+Dla8a58UqJFMRCDtj3OaPT6b6Y72d7dBQdW
KrbvGsrDkTum74ftdLXZLws7mJYS2D9jQKBMBfp2SlpjEAOHywydBEUpvj/D/i3yP5Xiiv17xq5+
EpRIRRlTZkGxlKUb0yaTVk0hXtC4IjKBjh+3HgtY1ZrzEggG+bomQ0ip/7AOZ3tm1JixXwrnADVb
uakhNubjy/IEUOO/MX0Vk3/QsREULWpQQXzkI3mWxs24shJ/ZJGBmcv5nd24jo/QSmPA+gEtUVIV
v3iPGvGGy4rb2QQhudn2guUICG3nIgAUeg6XzuEYsgks5bBcNbGX+Zz9A94TNamPzwZXx3bhh78D
K7VY48olRauSlz2pb+duqBpJcq+76F55KJbh5nRY7nWfZmmE0PdYLA6Adhz72PAE1NsBRhq6XEke
51Lpd6gTFsq93VZTBdp28bxjEtb2cKn+cp5vHN9hUBzkUM5+DlK1EaYMZa3Uqjm6KrlfOUWM981S
eX00RfIGDJqWe5Ex4X5hI+r+nK7YNWiMds1hM18yw8Au3Qw9f4Yfc7daBktTAh6vcVfjcNwXS+WM
pHV3f57D4BKZc3xa/xx57BEHedFuSFdBMBGPTQJhAOlEb+Ty5NLAVMgrdlPNXZ+gmGesSHenBQ0G
ID5b/K9Nppe6V4LJc8yfKXo+TSYYdCMZySh0fQp7pKuCdFviWg01lqvm912/OFYVhr6pzBE4BuKt
QqZFerIaLFtvS+r+oiQVaPG0O9z7v6BKwN9Um2DCZpz0OZ180P1W/A88mNHevxs9MGIE/k9b/otQ
XnlMvckNQ35oCXgDa8shIMdb2Sg1LCMo3XxtHEUYXACTLiz6gxWnb00At5k+/mxrTkkwH3ssJZXD
pzTtH2FtCaxlt+M3SIZWxiVYlKbNQjdql+zyRj9OCimOFDZT5c417cKveXEPxFTcTG6pRnZW67Yt
uV3D97n9suxfUfr0XDTGQlr7cd8sWEsegR3mYOOXb0RivcaLP/Oj3XTV+/spfhgm+Ibzd1AtQy+w
kO2xxQMW2MJQBx7FqhL1I9nPZcnGhsqw/rM7ONhWvo3NrKBeQYwyWwonucls4tVcoFTUgGA7MkCh
woa1dS0u5AhYRCcOQrjr72SQmlSoiBtynpEMChCuAOyKJ9q3en0cjPjtOKqepegJbIYCg2BLmRFl
8llbW6cCrPS37CmxyTMxWHVGTe2LwO1nJRZcBJG21HNfh7zi7O3FMJe+bP5ixdv9mtkzl3U1y0ve
0oPbSPyEkfjGg8+fKHbGYCAtrh8qu+7uLaXFVrdqEGiGMJf2em1oG9DgD/ILkgagGHAf1OX2bvan
Gdjs26EQzhqFPFb0Fcygiiu3nqHUjq/N/3M9hfyoBuub+WaD9iYmxoj8s7SX/oXOnBtAB75nWJ1r
KAobyqyWrUo2I7LJo4voOTsvxT5zI9sKc6AsSu4cjojJQwRy7Fr9vxGpUIGY9nvHAjTG98uSBBTZ
CDwuTrJFB55qvStO1vf6MRHSRGhO6Tj4Efm6r3IuEJVW1EsV1icwUoFMdosIf709+pJosk1BIX9P
2v/p+6ZU6mrDzS2atpbeJOhtyOvutwFBeCVs0a15hlHtWHJBiCqPeADwAaM7GjA14xqHb0hCW+f+
BP7LQ8P2Sz1ITucGS33R3Yl+IaycUx/5aDXzegocp+x47zkbjvjVAQi6txIoEW6SL0Kl4qZGxlnK
TwbTcR/w5Q0jAq3pPUyBpbBAfbqDgP2y/pgpZLF39TwufF5VCXsCwuWDbkb+Lzc9SecSMRdR2fXg
o8QeWj4QtJDOHOiRM5mVS2K3P8lxyrz3cg/S3CjE9WEkh6zCAVPXQqW9kXFsMSIobp49sS0Ba3dv
ef7DDX6PJVxAmV89/M61jWAn1/LuTpKRKljDTY2PMm7ulk/1GqmOinJc9o3U1AdC3LjW6e+5e876
xdnRY8wCuGlWoSat5cMgi1n9X8Fatq4yPJJe5b7rdVmdsmdtchKki/ec9ZWEwJNZm3j05XV95nEi
F/dsB499bF4dsQ1yrLLNzz3C4yZOZtZpGMmHZvFKjiZGo398cUdFpaPotA6dHV9AtJfgOLXiMQ9W
6uwkF8adgmsweWHpqOYeF48OmuGIRpQE7GoIKDCm0TRNiYF/4RUzGSoroBFR+dY7mhfX4DwmroFn
DmxZ8/GNv6GvTbh96/A5UUJHXdAzAmTSJrL7TPh9rbCz6ZjHkQ7x2TTtobw/46jmkK3kRYVLub9a
FuEz+/2Jhevf1ezRsis9oVbKICHXklnR5RuGM1EJx830vLcafI2l82Da2F013/7okJUDu+mPUto9
3zev6dXXWiDy9f6IDb33uWCb23n6A+nFFx3p2wWmZ6HtKHyRtjcykBGXcL6AU9BafT2nQOZvW8Tz
7zkWr11Wf6Og0J3bHNXQ2jIR5j8OrW+fBuNXCCsJPoDAeJ/KYj3PZqVoMXdDB4XZ528AfE7sMCtx
zMv8w0CtiOdqCakJxGQhxQSOkxBimICY0eireMGy5GZHmi/YnRZ1AXzZygmqUf7puJAr6Gjihj2F
5/gDA4TFgO0DLGjOAcLTD46KCyzag12/jK6iXHX8f69JMk9/W9EnFCKp6wBFdzDIezt0YPHjyUHY
jmeyo4mLUHqqruQPa1Ydes4+dlQxnAFRjnLgatFBsaCGGxVb3AGNcyUDAPoBQL2Bh2cFDFNGXb0/
tUl9+2zeLPqHEt2Gkk+UVYV8upUQbGq/FsjrpfyrvgXDEDr8b85Tpy2vQqo9aSSUCu2EoMnSSDh3
B49tOIbM6IMDW6bZw86jt8Zh03wZDfjWg30O660EAInWoxDTNutwnmJLVtlooQxpbGCRIk3aOC0U
WEAsMvRzYh+AgmXuuWF/YFVcaYeCuOA97gBn5n9RxLDopV+EOFVgnwmk6o4He1tr+3t3DjCQ+LBa
fu4ef7wkH4K+yS0N+78GbqWlhyrxY6d9HPZ/+mvcl9srTfcqavsqAUKbusMg2jDP9XaenNjo1trR
nB079QX8v7YZSAoKnlmnvHpCCiKFEzWYi5zDtIofJdUWnfyu7rvsKNWaYjJMuq5A2YrJIqHWA8cr
eSRx/llZOATWYsOtLwGGOY4VfyRcDBXe04qSDwzQnEPgoAtdFWpZG/jGU26hzvYndlKhkvpX3uym
mtBphPYIIn2h089ePifIjHLy9WK4mcT8weH/gOX9gcC5bTww4IH5f5C/vvMfVsnbyhl0ZvOtF56J
/w335v7z1vsYP+1w/WX4DgQKlv+watPnR3k8mg8TkV/1i/2hQlDRjTUJRSjzqrxbJnXEA55CtuCZ
rCNuweBflsFlJCaKhfQQNgHE9agnVEVYWfkaTRcXv7/2PS2oTVkguLIYhDL9pJ2Vu+virVOnSv9W
US6Etg+K2PJc2vPHPFIyje8aDwrZiL11zoRQ9mTytu4tgTP0Oa4yHZrS5QNpXOE4J1q4Ut4VOWAT
Wj3EOQJcn4EwSFBnffRzgcT/pWvpfm3gugj7f6PnyQPq+qe/UWYmzI8dISzgvG8N0weaMmyDtC11
FidKE84XIdFaNj2WQOLeuJpXALv0A6Hv8jpWG8A6bQYBnxWyUmH98uiILtmZz2nCIshnlDvntBoH
/ve9A8NOSAWyBet30l0ffv6M7tNLCIotV6mxj56jTOkKBy+LfLWG8dGbRyYe/jaGtnliz70Z/7+a
r192BJfY19P4yvL7cSEajEv2DFX0Ll75GjTxpCzU+/0pgQSot9dwn9sIwT5CMiJ5+5ApCT+dU9E3
GMtQcfSBrXVPJWGnTZg654zb3+YKoCvXNE5Eejg8I878ybiFMUusIQ7j8f1I699x2Hmq0ZHQbw+w
xjAcU7YmGvn2EBOgcfySv9ii7HriGU4S8S2ym25/kB9a1N0AQgPLlY5MUy11bhXeZtSlbu70LFc3
WYiG5ak5+lpssKCIsYmJCGxrdFWB/ySLaDxyPoHH5xIBdu8VgDh37brtkPinGieorwp2/tfgtyUr
QdQdctSSZSlA8XCVirkLziQcR07LIbCKfUerSDxuk6PrdJIiLidLZbDb5XEYucM0xyWtX1zqn19M
nbyCB3s8YqKjpxVs6HhLz5MU4GR6KdW6XUEAokro1v9mS54ba16c6JLTXm7DGviRHUXDLPrrZo4N
W7HuMmRpPIqb9ujXpmecHoXIWjn0Pov2ai3n2rdeXKLjBAbtwIyHjr4GWUOtvyoBRx1Ma21pJS2H
/fcn9C3jRgYbGzoYQNTjLpYQ7P5iMdQwKzmK60AqxeT7KDlvCiWqIIzG1E0S13TRCioshYxCQC/6
4iGgA8cfWChq4ozw932fRhKdGuUZ0ogsVn8A1zgwqg5JCggU6/0cVJWHLPPfHaB6RSayjv5qYhx9
Y6HjNZlwqf5HPNi7p7EW/Drl6zQifzHqLT39pIPMOZffevKj2ADzKSLLbzkrC0rmZ//l8XxCKCHL
YxtJIxCyacMsD79xKj6T7U86FL2enhWVno0n+n5LqNVbEc7dgNfQP3Vzp3a5IHKTJ1z556rav+nU
2iUdVUC/xqurekjczerNKp1eD5kCYuz0JCygemDifXILK6K5DEx4Xs2cJnCpJJS9447nYZirM2oV
7t6/8LAIKPQ8MwA22lGiBE3ErbgBKjMo/4OrJa1/NOw4GuJ/0MpV8PzAkuOtyeXnFYyafyw6q06w
kMVbjtzesVfT1fseXi8fZc25DO2IQGttS8mw9X4l+v3WkGc3a+tYHQ95QLg3wuWWv6FN+g5lbNdM
QFgLEGXpAiKyRC2W1eaLpR+X+5nSPNMPt5MLi7fYXNybQMQKNWqVsd4MF/bLiEsrT9LpFWl+G157
CES8qdd7Uzl+jTaMluK2zxNbcS70kqIk2/wEJhRYRwB4TEkfHeU2dhCU8N4+ykIN/eVGY2lKWXQV
SE7gUpH9HoMPX8rfRANRZL5mS24cXvXLR4wLfxETT79YIiq5b3kQG3wtL8aqDRYSmnD90/9MT7aS
xBdJuYf4fWb/fSuxI+CfUe6vnMpnxHw/w05Hs5z96MYHTRrz4DQD9aDIKhqWiAkx3G9XC8Z0uWnX
JW4P/+K0RIviV85jWgQwFv6To1YmWic8KKBSdo+VrAhH/tvPnYwrQa0JdMDPqaNnRbSfr89JUNcl
sfLzTwJJSWuO1SUZY1Gy3b0LY5RP6tRJLHwwzNULcD/nZqW/AHfme2uJywrOf4Vzop/IbQE9m1nT
MFZJpU6jTRlTYit7r6sPZiwEBgLwHVYs+iJ/7CEEdg6fDjrX8BzvNkkkJW0pbe4/kRbasS3I6htv
9q9IrW/fpqplXfjwRKgQ8SlWUdlY4uzDF+CtRDbaSHcNNDWpDpgTFUQvKcBKc3Hj8ZkCAuYLwwq4
omXSlrqcgu7ut6fvYXUGbTrk4HjBUl9iDPX3ow62d09UKxIcyFLhJ0XtfXUnR6RD0AwnV6pEjo1f
AYPgV1tHQy+I6Euca8nSArIN424QaVCu8V81uAWDIPLi4gRsxn3y3juNVLqzqyaslZmyb6BfjWeb
4ZhN0vAyHojHZNB6mtdDx489GXTiCk9D7BU6C+kMju9WVErQz40Mnb30Vl/So+bQ7bmC9GQ9CVSx
WqyOy9Gh0zUnwAzaeRzN02BMMADZWbVnb0nTwNFljHGZcgMaX52emiukhCA074mkCCYWNGK6egni
hn1ioICkp5qY2cIePRRjIMHHwLcJzgo/+I/jlGlzzA4HdHa4cfBR8iHjyU+214rGiG6GxvGkyL77
GloXOqFRbVdkRdcw9+o7BdEyKwqGAl2LtuHktVmrv1NPpgMLHHbhkZU8tXXYshw0YwqZ7EJqzz5V
YExNm+ab4bNDzSRYGT3elzFgAok9FiLaLiQ5wUV3/HItxRKvfEtaVafOM5lMgVo6v480B/Bvuw/Q
ezjgtE+K+D01RoCbBalmS5NZSbpviwfHND4HOg8DWt97yIRni5uNAaBnt47snOPGgDIxrMkOmm3b
U1rUuC683dcBvtatNysYdUdgF2f8TTuQe7VnTiRaDRvHdIkYq4yIWSDcWv3njbx9CpDSyWmDQCJj
/0utkrnsRDL8nv9QVIMkc52pTkVBDuZafhgOHmOu4fTKSBsg5p88LetBf+lf9GBQXalOcYUFGhAv
uuk9+/BvUl+sqRSnoWdfaDxsJLZYHGGiFCCIdINONsJ8NmVCfDtQNJhXO11KJ52PfUHConjYdGQJ
xsviZW3NJir6p0X2FuqpTEHjPaa8bDIKLTyBqtHhqxLRgs+hDEcHZS6Hk9sf1uZHHhO4T8hDOrG1
F4dJNTjxk/KrEZKJqjE7sxrvgVA9afwFywSkd2IEewowhLwNkbhiTYFZRQzQmViXXx3SyT7YSsbL
lRX2YOU4q3LHmNqJ9wOJkImaB3WhT/qWuGBZEVi03+JjTuj12bAn6620XZJq/4zrwAXNyU/hp5Sq
fhqwOv1FevIYELuQfWZ29Hb9PRHWJ++JmxnO+78sPw9z8O7ZaxCVfz3WFUSDZVji9euM29tD8xJ/
c1KWqpKHHwg3zf++rqimxELNwUsMaNJA64x1w2VeDJPdPptoa20/Lyuw99nQSEmOPYm+mdeA0E1a
TnQq2V9Z2ONKiMRkiQ4u62bqh77eWB9RkP01WWh5j0QGXeeiOgDRNOZra3YKNY+RXWVczGgcjfpg
7T/CYAkihXdAVzliBzb6qu0pSuz4hwNfGdkAkZoFMXuR+jIowaRsVPpwbSW9ea8XikyY9oDvrggx
nx5qnQe3N32rmCCJeVdu4evMBmO5PVPrKHQmCvVAANnLdWtj5pk0qWFaCzyZRZVEx4mWYEbaHjDz
7Sr0k45AutXr0XSunLooZG4MBXuAIcFUqlkVb66LC2J0FQhwZZToLPWlNJPWYs1Jq9dVodl2NVBI
MsyRQBqz4HXsiRMf/7M3Pf+6NfIBtz5B205ciBihCXcDB7xryMMBjCn50XQ97BSFzJqO8RdNvxKx
qGfWkgKVMPJ5kTtkQqYVJMSuEWR79BozK1x5u2ORGFp0xYjxgGNzKN0IeiBxEGCkQEflJomnRfiW
kiX7MlrM2pLLJF2W9UByx0jNOJ3stoaAtXM22PcFl2PM0mKyqyfQcpv5O2J+LjkAlsLI3CpKXLVV
LYeRbQ/B3sBiU50WgCZJDgRjXSt6sRbaQRog6LQkGJFDqvaim5g4aIoPpFEJpo3Eri4OIVB8mLzR
rreo2lHbVQIjGniT7ixYCwDdBp6QLEaxRSsrT03tDXMgP2xzKtT8hA48sxMJTQvveWR4HANvmAwa
Gno4v9NGSr1vG0PouFbIi1X6oOjm+ClxWESmcM83vl5xfN+XWmZVj/RgBdyaX4oqhch4EClwexc+
YRuxSIqAgTErzmiHkW5kMCJwxhJcDQAMruVygM1wEf4XJsQO/icNkFqTDww1W5FcZPpkNJ5/r+Yq
1BjK5eNv6NKawbLvtdNA90JuMPSO6iTzg8yPeHAcU6EZ3QavNIhWDb2SGUoWBSdu4B/QfllaIZJK
h+FhaAIMwNLSrlQyXVtq+Xq0FMEKNaRBcpcPHj/HIjnWE8/zo06KgJ5FT3j25qPDCTCxtZOP7SfW
1i2kdYVR0L3MXvxr2DGhpsa+sExXxy6EHo7hWPitRczumIszwIsQyy2j6d7RYHHjRjHPd7IB31a5
n0rkHFlwyo+F1V4UngXoFdhITVMuf2IaYHBJZ7YeIP+Zo5nAGfo8eCs9RvfyueOmdGUQ2tsTnvDH
eA6or8MdxIS0ReM4a09zW84cfY7QJw1UtwFnTc2bgRhety0tMtw7H6UhNkRMjyyudhWM6SXnEkrm
vAInUzLw9ioKZKnNiTQHTPy5HqZNvxx6YXAGFQU2r3Ha2YDwtCDxiJFoK836beVhkvR2PzEjimdG
jEuzK6w8Q5691wziyjIVWa3WNN2JzeTgNMmmvIEhPUcB8DjwNAyTu3AvfTekwMJwWmM7ORCvlql/
qzqQeocz0Hk7AbrVncoySPupwmBWMJzTesSu35ATkIakAPW/MC+n1MRHTqTVXHZvr7t+99mHXGR3
8bWhcyvwSYbdfOD6pORjLc+8RVe6S+u0Dtzcmv7zbtHWX+gyIIx1Sch7m5ay2C++QiuUTikycbfd
NC+xbIniIeoeiy/yt/dW5Y+OEHTSZrjHYrh3mS92jcQUaDxZj3Lyf7q8JdechA3UwWnxELikFwDx
4445uiNGtvJItdKmcQ4AcFyJCHLD7v15LGPAFZGu0X1Powe86yh9HXbAN2qs2lDFe6nkUYUOatV7
e6ViFw0qTi5vufa/LvkqoErTJIlrSHiSCd9z9CsUSUl3p7dw8cOuMbO/2vIccvdJMxjb73hGULaE
Bpovh8v8FaknIAncT0VWb8xxlLnaXedxPl44thV8CvVEdytlW6l1cWbSpgaoKUUxDL8ztjs4rf6q
DyJQUTJrbEBZe0Y04eaGPCl+g1B/YqKh6t4amjly6lISRfG7rVIs9Ls9apjj/uQuiB/rjC01Z8Gb
x9prMSTsHJQNPJravSLEw84Y7p7JX1nEOX+Y2wff8O6q47ayGMiA+zl/kBdEwK5R3O/D1mXu7BBv
mklm/1IxRSxJxmBIGpKntFozndAt23hmmWXZEtmB+dVKQdXp3vU8rYKHv6ql3p3N6/g1iWN8KxY4
nmCG+MrtNZgnLWbsUyUDJHmi4Pe/Qkt+Q8p5HuWgpcneXQLp9li1QBKEdlePUwl7dxyxZBuoZMwu
NDMnzqaEZp1L0O99i48QZmmzVD4qwvQJFv/wRd3/z155G9rAf13SpuYfhu/KMQqeM172WkBG+DOg
LQQeHGr7CT9jAe/VqZsTfzB0P0BTu6F8hS8R1Axr49glSwCx8ZxcIcNJ9DL7kbzDRxx9XkLnBgbl
dJ0zxullJqxInfoSgCswk0hA0XUxYlk7PsVNYiVt0erZxzNv2Gusz5eEgVjTuyuPNUf/JOC3B0Ae
63iEu04xCJKcfvaKwGbSIpiISun/OQ/YiKFKvn+MIyGmW6jZPwt9bkahXBIwwdNYoDsOUuGbGzYM
Pbj7srkc3w0M704PFmqZvR0YejXtNDsUjoK2SgLrShl/fSnQqzt63YGqI2UvZTqw26/H4n8oEkEs
OYEmisc+g52CCJNllhMcY01IxUyJm1q80CxHWBtzAOJbW8Anyw8TgQLPd4UJ1BwSp4dSHvSYZpvV
UvIN0MwcgQKbujTiyUIOgBB9fMdqDt+lv8WH2sfsG8bi1OHuHDqkwVuQ+9j1whAFrdayA9fQ8Zvl
HoYK/LSYPBCv5VuedNlM0dPo8VM+8qqREikuEYpo0NvR7w9VamsC0gB3uUEHrO5l4zzFtKi8ujRr
opgHMdi5Cq+4j//qNDgXD6jJFHJh3y2zzwoMIhv65L55DNN3WJZ8l6+6rpZ3W+MF0GvY/E+xom5s
kV4QG1x3bLlwENuEFZv2SicBqWxJtPwH+Z00Vgb2W61lqajzqay4aranEbdWp/2nJO+haX+ieJay
RBDe60PQP8JU08Q5+2p0CW/3BhmocX/epX1JMOSb8pphJoYyLXlkU9EIFbG9E5tAshRmEg7l9giA
g6Th3yHl5bFvh6jA1OPDSjDrO/xYf+fMzqEtrMoDyryAQbaoCPuWgTTsDu/Q8/yY78sETX0X6xUs
YTxZpW6CAHbhAblNA1oLkTgKwpJRrv3MRD0y9C4HiPifDnbiEnB4COB2F7dNkqB72/f+915/Axid
RNZNUZYKQyLb84Hu/c5ooSIqYhzmVpx6kiC2ygb5JZ27qUfn1sme5A8k1gD4BBEOBFMCwlojbdnf
6CYctZwA2P6TxyKwoe81ekLD/MRzeCYc0iTEakOhg49ZQYZLexOwufAsazUk5RSqbtvSamNdtlAn
pLVPjUBQy6bzaAjlmjdn0uqDbAsNv4tUFGh1DWdQ+xqstv7+D/ghRj7p1cBAo/DQwFK76VparoxX
yg2N64rQdDra/okjq07ky7pwSIoZLlwARHT912gFH615sVgDi54SFrhSGqq7nEkO88TqFn77VTGB
Kom8JV9LqB/NVVfjPS1Piba660wSsPEKs8RWqGzYIZ4XRJjx5Utc7tuYdVv07B27YIaLmKkftQs7
sIY0X4u/vCtSyyNd7Klrrfjp4AKWS+R3P6umC/9j4cH1bXD26j8vYED6XCuWuMh+hpoG1Z5I4de7
3y8QsiQSine2VnmyrYHEkIzqiwu9jVUiuuC78yCpPhaju/qFP8uiSRdJrt5DaXVzfaYtF2fVIOaK
hsLre3x2qoC2hjMtBimzZlJvffOqQkDyOEeIoB+4kjN7JiTjmjhtr4e6NHVVx2FC4IKev9vQMXVg
+gbA04IKDDsFGmJLGJ3cp1bBkaDof4VGrRNoV6lAO70EDC1jW8nt/MQyKBj+l48sUXYIqMneAMSV
dGjNPf5F/f1LKH/2soRH+DhueJ8qSrLRlwSrhSjL6nuHt18hXwW4cbie3xGmHNzKGq1QNUoyKw+6
oQ5iKtNe6q5xL0xawGOTZh5hMawXTCuOMlzDg3mW+1CE82svcRX4B5Ds6AZ1iF2BAAL7Z736s7Ql
ifZElmYjUl2vcbyCcwkdqR6LrpH3ez2bRxzNA5k6p4Ewwx5hmlbw0ffc94QSAy5C3cX2CAdXyKag
C8ePnGwdwGYj15XgAteRKs8POamtiWVVpo0sPWxIycMR7nKRzErTAFwFggsWn2ex0yNzZK/t1Tof
molIrIQhQYLWMijwyjbRJEDfIeRRTEqY5no6Vf2DwMYrn8Gcp15whT05QO8VEkCRhgFdyaiUU2Kq
+GcpPOWDHt9eFrQqF53Ip0fXHriw5tWeAEP3QfYUT9G4kJ68LYNBhc4JcQljhA5UwiDNU4AiSlT8
CUu29FsJkeIiGRhfgM+pZWnqNap3U7q9WDGNsqOPpn55yE2MEOZpHlfHwtxbZquiFUi5yONOuXPp
RMq1B+uGohjJufQRQUbArTQOJdHSQOpqOZkuYmBlduGl+cYnereDvvHCxIclqW27V+iA4HNWt7Je
CTRxCsEFo/cQ3lEylKufBfF629T43Y8fiHh/AbL6fjb8VPozitamR8tjaZQn6EpqGY9lWdSIoD8y
wYaCfoOqmziV0ofKRudCHSpo35VCQvrXEHutu+FaGFdkp+xiMWRtXu6pg32Teh949B1eKArXvBfv
gNVZfF/OY2wSTdOG1oOQJEki1Rp9FQ8fVJ1u3zQxFKT2D59qXwSsYdAszQvf0acYQUhG8YHQxSgG
fZWgyn79AyXpmF0OfObJQfT5tcJDF0gnT6mJAY7L0bK0/y9s48exe5yrVEeD+BxdZtXNipE/eav+
AuEhuy/MCHN8clDrdVsSKU2D1VrIy7H/qOvk10PegkQPQHTeWSJltk1LhdLd8kFVaG/QIBnmRklm
8WrCHFG2ayFfGV1fMeV097RvQKTPq9z541BWcqWMK964MnoBOP/QJFevDCe16o/162RJiR4q1qLU
fl7QhEZZyRWQqrTcysjhrirWWLmVqkL1EO/fOI1RHPNFy9Aw1l+4bHJzhcOabxSGI6YmrzBqvcQ8
l6FChr5OUrm6thEyQB7OLYx2MZh1LCk6cMBjSOyK06FDcuoysITmb9Rysh3+6VXKZK14eXJ3kdcq
3HRB4qwJrc0YeuIyxOjoUdWsm9HYAZPzNHC+BN5z5wtBKUdxLZ49h2DYoB+9rUZTRgmsXnsWxrCx
BwU/Nr6KFq6LBrKjPT8Ez2ZQlYoJsz+fruShFq92q8ohOlO37it7rtnTTocvDJARobxj8oYgoVO6
mpajvJ4cRDpBn/Fl8zfxf1x69dQodEjBdNs/zm2VlgfgHLihwFEJnujXuulC3OraHQf/RxWNo+qR
oE9jCsdwrY0e6ThZJ6iW/g64rNtWzGRqLK2UBe9lSWoX3agxDDUbKA2eO/MAQMgIOReEFmVQNdSf
QCuxkqjy5LA0ZFKmcJIhu8WK1rpbW6LGu+5fvE4xoDOfmxX4X6ZmwsTLyF7HrgzMD0ojeJiEBTMC
TqdO9amvB0YEjG/8Ci9Ne2CI4+zGfcQEQCjzHfzGuIl3giSl4Sq0AZC5/u+U6jht6UcAIrgAOJAf
w4q4/8TqXic9B11Pxql2oZFDwl/h7Y9vN/04U6tWiErahfln+QOWPVSpQRgti85u1hcED4WMZ91Z
KvXE+BufWGcxCKQF9uiHwmHTk8fF1FNLwPQPHj0BgKmcNmWEser0ipQNFHaUNfT39SC+APPgg7lV
5dfza9Ng+mU44dwazCjrJ7OqdiJorrX0ySeMzFet6sSCiCH9ZFSduigni7Ed2pnwycv5Ms3MF8hj
dY3S4YDJ/U0TYQjzjRmq9riBk5llyQb7bnReXFdAR/9Ulcs1xncis52+4SDWt6chJ54YhblF4TQE
hYtCPjwxbbjpE9fLNqtPEkJTi0QCePTB94os0TBHu/u7NoK0jXJTV4fgyu2qHke16LLaAeDgEuNc
llIzBCDirz2VVHdtYIigv3wYcUgxuj54ylFeZFNjgHWzmZS3kz5yfsuByRvxh96poUV9wJYfsHi6
qgOzIVXkIUwr73h2swk0e5Ddyh7BjK/kMA/wcd44Qpg0BnUJHItTXtvlUibQ7OLcQvCrbXb90y2o
QdcsuIDxOIPXl9pNnwRG6wWnFDPzMcf15ms4YjkRGI8wZaAvc7f/4sWnUn15SabBJx8vYbITb5Nn
JpowQPCwOV5R/uR2kZA9zjOsmpSgVDXleD7rSlqsj8ZhAUJTlgNqOpbq//3LvRaQ4g/6/4KUNTo+
oNO5giHg/ai/Tjm7Ey2kE7MrMUzfvPoykOC/x3E4ct5ao89iANNbXs1Bfk1axUqZL8f/6uVRVrby
WtBgnDR2SyjEU4Pm4+1Io7DVQBm4nJKp3lHqK+/SZYt9r2ns4OG6LwP5DjKleH6GZ4dL7d8O2b4q
9CqRM5vtqjpOnM+K0ksHP2+CLHrlPo1IerWCd7ReBOvyQFBZKlyy3ARtqBzkPO/Q0FeyZn6IjTYh
p2IRGtGNJHQ8Z/E6NCqbBs+atSujryFD0VpruSiL2rS9yu41xx+i+Vih8JuoBTHL+yjlcEttMDrG
BA0HojP74qadOF3EbTSCNRFfHxXt5bQYhyDEHzJQBefqul7usvyOB3o7byxN/fuDjLWEEW3LPY7N
/+h3CrknqB7mU0wmFpYZntPaVFzyd6NlfTwVwU21M3kREZM8VhzaW8bSwUrluMXlbXXY8S8VCae4
0et2OPNqvehjYHwworMjOnPZpng0e3/7vi/yjA2+FlKj5Dje33CGdD96D6i5kvKNbFCcI37otpIJ
U+Ns7Gm4XcUDMHutBYFTXJpl34q7wJ1j9dgd43oCW/Eg1S5MmnurEJ3uwCMD8YWA8qTSNhZOOztv
Y96O02oEcbiWPqnaZuPwUsd7CrceodJUBweX7XPqBF7Iqt3iJBdXo3YhaJXA0l/RJcI/uQSBqN9o
qj00gc83V2g4IL9ovAh6vsRt8teP+kmerOKsrqOIUbYB63SANUHKDg2K7/ZA6IHbAZe7JG3S5E8F
qSAwo+vwXXofFyFEjorXgUEswogrY64M6EHkzAWmqpghCUHw+tjuZbZtaIiMPfanvoOBXBJv6z5M
WUsgzb4Xv4fm45FO4lf1Y0hb+G0P8v69A1NTiCDufvnWa+C5zjn9Jx2wn08IwSIyS5qmD7zPiOG2
BD1sIQftBxmy99q0qyA7yDyHj/5NwSU8equ2GmS99gX0oqFV4diB/OrQQ5qVJzpCTwF6ql0tNa2W
iqYs9MaYvAhToiz+1iYL0Z1rxJZSaPQ5M5KBL1LFUaUrlZ4kn25i+YP2AiaG6gBffks3FxweNlLZ
Wjekhgc3gsjB3HTJD+P3nCxUIg7Z1icMOGWhaSWIF224eYWNRH38qV2IZfZ2zkRMqM4B4AFW/drv
u5POojK0t0UlM6El1ghE4tTa/XRG9JbPQN3jzuJkidXuQNPx0rQpQhdNZ3xUTykzAvS56GvKRB2z
I2qz1oHbTV+rjDjPGK7KGiiJQbA1rcgUN7mXdncdxpUDOdNfS80mDVAbc7MkZAeGcLihV/sY50YX
FRJ4SNpng8l9ffizZRsBuCfcMWQfDtEPHxMd/X8bR5qizaeR2KtU9RXS0hIH3aF/WyGs69kmC1dI
QDf+qIYMleeWrR4e2oWTcNdcty8pbTFiOnVC7Ukn4xo2X4VaHJlNJbYZi5UTAD1kegzmML52hKi6
O/rj19pFIsP4zJRLWllTYPg2RLC3xH8fPGB9N3jA2wNpOxdbuFPs8n4GsBasX7VcP1qcDtnoB9Xr
LtUEhmy+uz6BP8cGbD4bYfRZ+0uLgIdylITIcRvBqRMW6BxHIHo16+yS/DlZIg9qWOllAm4fXCRF
VlW1kIHhl2Jz31EiSUeflUFUjd0CYV7o3Bc+HxLtEoJ7uGOFJN+ovHkU0naHCvglrTaZcT61qXED
ncGQWJ+Ufu59jMwXLptlvHWDad1wBzDfGwAUqNkxigF43rhPGqubAh5ada+Vvx9g3ys2iApOaLzq
JQeN1a5G4KwAzImRtCUayiEZeejN8avsBd781q4Na1UkqOz+sCC5s0xS6O4kaDYauTWfGUIGfL1A
fNiVN02DGRmWbSKyWdY9BbCMTA/+wfFetGmfkOlpnQBW/mhpGjNs86lqaIO3PNatploFcWaGQFFx
niZmYeAhobDxI1CIjo5MxLjbfXKJiMah29m0xO6H3lcb28Bb/uHx68VK9NqBQk7eyiDf3uI6mzo9
VQOCwYtCYupJAAY2Bowt2wl+AxvwfR3RL289pFm7r6OupwZ2L0zPF1SQqOmL6IcGHQlBUr4G077b
qW6qz69tdNdApaZwjtKFYXJtwXcmCQDECR0t8T7CXR7iY9hDCrh+5o/y0umYy+2df40DOeseIbKE
Jl8j2CMTuW9mQ2lo6Y1ETX+Y0AupMkqxWTBwQuldpY12bjt/4RDQn5K484cgGkzkymQdzwH7ND3A
Ui1NzhkO3weEz81//BwlLaenYgRrbxI5jkEoCEZXiTQeQKGBK5wX6qjmc9+ZUcz+Y6bgYNHaBStF
tv8LzAK6xs+I+hqh6Gy8CC6nm7xvWsDNMpqMW04qyr/owt1wwnD0npvvuht2AZgE6hr2F1Bdn2Qg
yHOhp3gqEehZRrLFH7jqtHa8CKxoIIoeQjyx2c8e0nguT4/3Pp1JFnnraAkh4LAF44rJHXB6F+ZK
5DCQa4RANVw6bOs+Tt3q0GQWjVAfZcSeoI3C0ysIRbBi/O0r7/Hiq5Q/c1WbJ4AKQISzj9rb8RE8
GgtaBRkXQ4L9IDcH3qVDULC2/DNBmZFnyWZwHscaWLLtH96MM2ONyfEzBtp9rj1rhD/uejTRghm5
fTj6lB02lYn+F0z4rDcDBIspF1wUPsBrisvjBk9FUR1T/kEN3RymsTEU8PQURYK9tzOWoQk0f7Tx
CAaAoNVE2fiFPFRdCJIKUrGwuSKnCa9tYlY26Bv5i01mH5rDUR6w9czL5XwdHILctR3BVU/M9yGZ
yjXWOZ/0uPoCDMgUFJWNnJYufvcMM0DPwbqWMKpRYX9JZnHEeDuyz/UlnGvK107P4JGJVxn3osbW
Q8uuVhTm12QHyi3E2Ybe5GDCDrgToppSbfw7iPpzEVbmdyIXbAhVQLOfUygzoAzkEctxQA6SWp+R
5H2MTgb6KLSa9CHVG9iHB5u+CgYiWnnBx0jrh6jeO7fxE86P/IjXBYSWYPSG9BJ1mT+ntaAMqNyp
pB/3Plcg9+1G8A7EWCbWC7AZDMz+0WChdQtFNTTraRSK5Esu1l8mEUXqodz3wtq6MYnWOSwXNzu5
KnLtPuCMEFxCpZTrVJ+i1LuNLFIeWRRG+bV0fTnMwBfdyMdO89PL1OFAOFnfWlF8DuBbbWia7p8o
IGyerORKcLI2UcumVcpn6mMmlZi9/JejS9lErahDVAfaU9VS5VzOCBX/dXWzGp5RaAYUe+0eAbEt
cCnDGCQuU8577EWZZuBTNmHt9TVNdcrgDAaS2cQJw8Rby5Ld4nv/gnlIW7GMdT5ZY5KxORZ404jk
fuJYCpMdkmFgzxX2WenBToAvgygzuBYZu/Spig/BrZ5g9OCUvbDBLQgYMrjAzSUFYbKRjmW0SgF5
0iVQPqG9UrXL4Ebg8VDNZtRlZDzgHIp1AThTCRFC/LNcErWKg133USG/TGhJlOtkvbO0ItyOVqYx
KrNjktMu4H5cOO547KTKQB9uuCF9QZMXGf4vyTUTlX9IT3o+Z6a6ca0QAiwuvHw4PATIcJVARvB+
hsRmmRXNLlkTZOcS00x7rCrK6ICFZ3Gwphuwxnap5MbTdIyFPhYYZSiAIbM0XbGl5FRJDmdzdper
j4KLpK+3K+lnTT5uQssHkZ535vnQU2aQvgNBwRc+Ycga7AOwLcMQ27a7ewSQ5AjrRpw2YItqhbfu
lywyNtuRBHStR+J0oXz7e8Hmmmrc1PuW24rgUkAPAcHmToB0yRzEhfMOFMajGWdcqTjWi6BbziEV
ojj8ZbaQSIliA3SthI5LyLIyeUHprg/cwsTmSw+DLGzaOcrDUlYx+TQdXvjDF7QZtMHeTV6KvLOr
JTATdt3OorLLDuJGg04Yi8ORfRTj/GqM1dEslRiviWgob4DOiUZPg8TvqLQKJh0SMbh/qKwVT80P
HW1r7yhkrocsj4OIcytHZHHm0911IB9G3K4Pn3CH5gwNjEJF2wPpQioOfNo8MY2MQylLy5uqFQsT
Cnd8zo7sUZtsP96PpwlzDgEGZ963SxjL0cR2t5/GKsOHC2BBCemfc5hI4bEiRzEP1j9uIkx5o41w
xmhuvtcpRIBhDEOfKPxJEctWm5nuzYrxebo/zef6kEo7/FGXF4g5ly5Bzp8fBzxqP+Kddf1ifAsN
hAUtkVXKR7rhbSuB7CaUqtYzQHbFKFBuqOi/W41Mn179bMam7agWedXpFDinPb9ZYF93qH1X9bzc
S+XBpcrkbkwQU+FjtrUOvQ7xkg/Am9YPMzFeCoeMMHcwc+kJvuZBM1pcl+cZSbNOU+/+g/fC+h7I
2NlX3upsnh9eCOwy2q5hvpK0W/cRKdDu46zZi7Bjcz3sL8IPj5XwOp8UlT9+SH6dmw87WU93tPgC
MwyioEGODpXreNTzT2d2aNakNRetPg36XTNuNl0dDE0SUNmlbXbY076mDgh2BB++2AwDOS85Qz1P
l3q8ElYZFIuPjdE6XulGdqJsXI/ehaOwsMokKaCXD3SAc1bHl+JyBi97I7M9fCq0It7YyWiUhwoU
o4AvbUtunflEhucAeQ0Kjj6sua6bbE+FTf4Xsf3DwseDG0j70UR3CQcXgvj0FpltqlJhCJke1dH9
dXo76WCASExV1TQOooKuPpjCA7CSYaOsYKD7jUq1hv1JnwKDo7EKbKk28T7iSFb2FAje/wIaOmIL
6wr2RWVtdNL980qTSe0YnA1doWVh4lfT1QWUKTz7uScZXEQE8r6WYwMCuO6bEGxiy6HpV8l+0dRD
MSzBSDliKN1/XePjUIAr397mXWVoWPDtZWD0HxGVkVZ+2M4PgzJXzf/ev44OkOwOUCpjvB8uN2Cw
R9LUWJjuHas1nz/J12S75LALBjx3SXAVfnDUlBtFO5e8K/5Zjk4R831qlYVZ5FqK1w5bfkSCHe83
3eP729ySeHbTl5B4EMlyxSrHOi8cgKt2S8+M+unatFMJ3VA0DovLjL8AKe9BF+VBFKh3wb+EncwI
gQsCOe7sCLA1bzzhXE/IeqDJjB7BCpFQ0PuqI3+NgLDWqZnQh3St4zIn8LTLI9nABb08pWBLd8vE
AxD/GwgOPmSCnMa1DEjFTe63mKfRAZkay6UnEU2zyPW2cWpMCxz3sfpi+Y5kK1QkzoLRFBXDwkYw
zz76WQaffAKrHgLnK6AKIoFkOmsoDqVZ0PgBofeOF2NS8ONnTZVy6hpN6f4kb5V+RaHI6jeBXEgl
rcfgR8dMO5K9Q1tiaibLQmuZA8J1v+0vA6LSLMdGLz3/d18Rt4/6uwiZlMVp4COTdOF+0OgDTQ4L
UZ8K7OX5L3jH/e/b8mD31Hk7b+P4qU4XiH31KTWtWMV+JILCBj2wm8M+tVoAOZXLurDdQMW8ap9L
CkqO0Sigq041XBqTsz0bTls6JwyTLqKo+RPAymKcmoqULzoukoY9zR8eSVpovmG9B+zsmy1HWm/U
d4onxnH9CGffIFIlFuw9tCihHzee2ZQiRhxf8BEmkcSo88wkn+zkDD3WfPIkLS+rWyFqXGjjEhe8
27fiqn5mxSmkfceG2YzTkQaqf4U83egBKzmemhp2UBeeM2xhPsdFGK8266vLExccyQozC1frpLTw
A+qaHIaJYeEKxG6kGlnOKaItKyt8swS1KO+XZ956IRA832VgYHNhpFc8e151RBnTx0IvSdRLPFWE
WKVssVcSf93yT3OAfAhTtaqjpHlMSbO0NAjyeHvDhtfX8/b4vUtE14RJsKPZH1A5gNX6QgingW0Z
dGeqvR1e99b5JKjbkAtJ/y/eXK+r3T7FPWhjGCqMKzvyS/p343BKC5Dyx1sEzSJrGCji/woVQ4qt
25/yqYaFv+QEqFmPMJtr3HcscofHRJlhR0VD6ehBQN20M0j6y4zf01nf8Jlb5/BiNrlSJZyzicaE
Q27oj9I1twx99cjQXN9hdNcFJCBKF7HQgoFIagXKZdWFzWqPwt0I834x5Wz/yW3K5UeBUxo/zcMI
rH18RHGr1W6efVx4q7x2+S8VaXIH3v2L6M6xjXblqr29hrxyMXUvG/dyOnzRcupYRQZOdn94Yutn
XUK0Q3y8RN6m6wvrX1ka9nMq5pEz8Un3auXnkFtB9Q+maof5bhBJvNQ9RtPiZjO8dAmie5kgiVwC
XpSX8Rw3VzMezNXymX14OeInfmTpfvSK1jGa4s2+P3sa6REjwMu4Q8JUmuz6GsZRPWmUCz/LwPLL
NGIxc5PbPXFPAaFtdR8p/qybj5rYSeoAeKWlGY4UguXBZn7cUkmEMBQX13pPPHXICTOTPD0sI5zF
rQNqWBMHotZssWRcqpopisopLY4JJPKSv2lwhuUs3s3k/SN54o8jjxr+xPQl/SzkIIyMnFUhx0L8
TWN5GGvAos/6pRKNpzBVoEps8rLkFR3EGV0h2LgH63SiXC0eD0dfBhoDGbzdfIUhy4865a00c3HK
cLYEo7zVsq0U5UL1ltp58l1feMWANFzzu2NWCAx8foZW5UdVKUrk/rbr+kaGTV0ZG3zHQ5rMRyQt
znPiSX4HvpQzGoX7yhnc2a3jh3RIaeUIxumQFQRFHVQgN336Qkd2fsXAxEGkmVpBiMLGc8mVMYb9
o2O4HpJaIJFxJmiR8+DXrG7Lvj73mi0Ws2/KJrytl0QNeilNo+bPUtpts2QFIhj6pXxhsFRDUywv
oHKxyd/Gfyk3HvUKuUuWZoG7fGkR36m+Kig6QCSojei5iAKlqw1/REiup3ktAoR7LzTJlweMMig5
Dr1UhXJhZPzB7XO43zoH1GwBOlZXfpKAov+LR3BL767xKLBJjk4L842+I4N8ngdmmgEOaHWlXBzH
PXm8m+emfBYpHjJc8X2dGrlE64jOS+SWB01nK/ucrNfEbE9YD2yOOxpjGAN388PY9YyBMesHGlfn
x/Pv41SMuWdZtWwKGGSwLDeSUN0P1Mmc2uU3iBuUHgO1ZV+63WW1Qw7VvsmJxKQ6tPNiT46LmKwO
+LNJ/f2POulOWZDSlzWYVgu6v+QGM0+ffchz86674i+V2Ma6nF/FfMw6X0QW5pLc0N2jdGFePFV/
YvxfUmuutGqbzvZAk+LKRGv3ZvE8oGCkl3/i6fpNuOSbyRQxbelZygdFEEJonlYG3MhK8CmCeVRd
6A6tEJC6OFr0epSlIgZ0/lHJGhy0SP1P3t/u+d+0fF96j06nDIAHbJis7r8LmR8TucZQ3ylJ1tmX
bCsIjkmyOKZYJC/nPRDgpQ13Pr7UNHlfjzgkdI1pXl5MFzIBn0KhawV8DaZLesWmnBNfaiCSsbGt
wS7TM7Dsy+mLkBRh07FGKLts8y2M81CGIAU87oVyt+yUBBVk+jQPA2AmoPcocflJGaEHc/TuHtVC
M2xuS6o0g/GJuA4vllF4V9LPFKvB+ioeyC8DOP8hphxG59ZPRiLxUXJUv0C2pU9BYDwl/qrFqX/I
J2gTCNLGg3fM5mWTlUeh9wiZWOnWVVN7zCYyOQv8bGxxKEYAsg9FQBmhMiuH7sbLROUGnNYuz+dd
RmO+ITES7AHTZtb2G9qQxk7DmMdnhJFyb63767tFJ00ZKm3xE990njrB3lF/xwg1uI5r+CN+4Vqg
kEhkr1JVS1BReK6AKTeDkDbEpvNB0CN8h1e/awLU8mWkiqUMCse+6fe2wb8G/ZAw4Xd4pLD+qoq8
rjPsoLR0y1fl/yv2a7DEQhP2JYDkdG8JAXsBMFc1z/jenyVtv/YpNQ9FY6HgsguXFWwfp5hCHsDf
lNvJQ1JH+LKZ2PDI0kmgQyC3gLfT7iLXpmQocYpDBUoonCejliVJstsC2okoyGE+eTo7n94kxoJ+
PELJpIvdF1+qVldqj7as5KN0CdHBjUpamqG7fLay6gvdmTMmQOfuD4wLVDk4WORsaZTn1mCDgCB0
9AjBRHKKfhRCqh9+KI8wcBtzGhc6Jajg8jmXgz9rRqon3WXNkviubfd3KQYD81t82onGnVb9Grh4
8AK8wFzFILzuB1raZJyxITBxHRrm4NcrnxPIYydxV6/Fqnp4WaAxHeGU1SzHK31nCqI5UYkz0k26
lBzoV6ICNBaM6kaxQIGy1jpTkO38Kz08JEj/ta71k0wXTSjxwbxGVy8235Y8aVTKqikqFtB9kAs1
GaF/S/xIryFXjExZqkYj+kuLXNbDJrUvKTxLXnwXx8shbb1613d4D53hbmKQxOix/P+v4EoVrdYA
4kYg6FXfSUUd98sroBUOQ038fussoRS86e9KjsDzvwTXF524cWq27VLyU0kcdlU+t+fcEHwxZzB3
9df/c8LB4hX0aqazEj0yPI8cpbf3TG2m5pSx5BRRoJE2o6lOrMBOBk/Ab8fFTeXaCvNbNJ9MDzk8
h5SnUi1UhWLMBOIRcTYFR6XknLkCbaxmTPgYhSjSZTpYPSnCdPLKuikFk7134xtcUODgndJ2qqCH
Hefv1d+X+QfqfwpcXMeJ0VInh+vF6aT0sth8cncrrHemtN+YwWFFY0bEwuxTHiPTlopwEkbMCdMj
5nkasQuxIG1b92hZCQDrL6eB6lnQXSD0cvxMsNAeJRDMPHggWaG5NLZy6CIKCwP9ntCgf+hUcnxz
XpEZolqwVNgKKFZ0vaiKnchZDh5Z+txCSEdLEi9VaKIVdbVtasASXN9p1OBVSckO+K1omWdcw8oS
Jl2+jLaR2gzuhr7LBvE92cV7C9CGUux/+i72qwItfa4hRyWe1YCDGnrKgxtj0i2kqYtnUcEh65Xy
bJcFvBOwBIEJmW5FKRg4t+g6hF007CVsQgAZO9ntEXAg0fYFtZ919kst8lyxDerSLG8xq83PKduH
2BKkCpa1vR85jMlIgGtR2MJa+QTak0p0H5wXhULPswFDanHsoNn8yT9zT2q4ik1k9oKPYg+NJjyM
jTbZMQoCv//POn1bL1pRFrM888v/XRok9w1o6whcPoo5923cdhxsd9j714o9ri4s3bYQV0hoOshe
fQqfRKoGPSK97ojqQlvPeWDfXmIxFhtHeIB2m9U7Gfndjcw1sI7TjbOg/8rM5qXdJ6wxQA7lNgxh
XPgpIwYK6n+J5I1ZEUu4v+Kk9cNU4MDeQjxMOMtKhdMlSeNuPhmdxSsL3EbcLzhP/lYm5QrAdDdr
HYhIUch816+MB6wybPA9sQj6kUFZ8e5fQzlXs1snYBfrGOj23t6zS9pWglrhmFiqSa10AHg9hnKI
8UBkxxPmJkIld1buRyXr81t27LnwOJ4tLWci2rpx6uGCKCqVd/V3xtOGMN6cDribRkKF5pkzj8e8
jTtkoaOq4CoSrcth5DEuSw+oCCl0jelqokaV3A/Vy96yUYbhKuRTxNWOuDbH/R2rC7SIGxNkcyaG
FSzBlugjaKUULArZYASV2Bu/uXLOIu9OGNyRefk9mp/9vXDsa6UStEA7gdprOpC42UsBX5R8ROeE
4R+GC5zYFuUHtBhWcBIUKbnMmSZ8LlZw+ALysy433omPMRUKw+jscrXCCr21foXX/1HIhSiOvNti
AffRJaNmdI4ChpL79sm3CDbftBdBH93DcJF+qH5w9CrlidPpX/KSmagVkN4WXuaCFMdjN4tzdalM
dEO/wHwK8wjImcEZZiBTBIwoa9JoLh7Il6twQzfXyxyd1wxdqNOmMIImlvuQpDEgV5LnX1Zj3NJ5
PYjB7VrW7PB84HpUXk9ahMgowZDW/cwgRr1hdfOLT0n6tX9/8exLhHMtzs9UaqpCcSDJPLDYtb+n
B8865kh4PeOLJLw7qTVpE+FK+GQeCG7Lu5I0juflBMjhlHoGDswN1XC7qFjEIIoXd4fbbSlWPjb3
2HZkgs2MBHyuEVvGVrVbAnHTeW9KeAbsSwoY+dexIZ5AHxB/4B0npCp8RRAPR3OjHPiQ4MmAaHIO
5XcMgKO/nkSs7Nhk9qOvyi0ij/PxSjOm7u6Dw5QhFL12jHsmF5rqo0dnybMp0K+iOxmP6DAHopKk
ZrEYzzzhv2Let3ExkkXl/GWjx7SQlcrQQSCObRfe8ujBkb9YXjXVtK1PD/GNf0K78RcCuDAOb/+K
1Do96tW1qUtHhH6OdX9RIxigzGLMjxyNJZn9zSU+g8KbEWZ4vdLr282rOfxxNzOla7KfFHVbolq4
QJR8tbaXdRulXlBExxToF/xjjlBhb9AuffSOnrvGYOjaD7XLoAb4sLLohorV1F0dWfQMqe4HLIjY
znA5LUzT1O8w/hUUX38qXNvGrV+8lh5c9e1hTBlpS2Iiymb7YP2NwuZ049mlFMTuPZDCibR86CKm
ii/mQTKqipN9mrgziAcrrz07YEcuB9VzNDJothhIfE8VeTzFH1Ilqkai+351rU+zFFPp/e9mCz9p
UP9YTiF7wj/inKS5dn8eRb1EcEW7Z0MqB3J63JugQC40p+DXvAV3+F+UIh2Zq1t2uOqwNcJvtrQJ
tOOUnif7E7Pm/pjgigU00jAlka6PgQU3ZlDTVzlZSCkixFb4Gv6HKpuRVn5ENkXm+ZFTB99thO6O
6ckRBUtPXp7YxMSVHuGQ94zcN65dQ38kFnssZw+VF7yAeKKH1Esfn7kaHa0+o1bbpsjpShYmtM0q
TzLWLMH2E++AkUAlI0SCsf2XypL5g+hqDvFV5XufiBv8FH2lh25o1wXp1OcFIAq/1gs2UxdVDXH0
Pn7lzoVjUe6dEwTUsWyUlCDNW3dgcxxGDNsudKntYecOraY6eau0bxcjv81WpDWufjkNJ9VP9tMS
68GeiDjhZpiHLFjiRrQaMIimkslRTpcApbhcsZguIZ1ht5E7aGDytjgLaCFFbGammhaaiRZu7olJ
an6DbaoQ1IRNhSa0UOUwkF/ajPBro/K4a9tpUcdVkP0pZXJ5CLj7sc1UZS8r0Nj6QsG6zFz6xB0x
42sUkd1S91m3HfwTpi5TiaCgZKSPIHpzkBQkQV79Lrb4Bzp1NUgW2ASk6Q2Tp6q2Jve82IXmaa2f
BFTiSf+ilnlu/X1ov98piXkFfQIMSnESJgCnZ67pqq93RapevnsbkqGW6+gTP7e+vp0W/rjHjG3I
mYEJIiFkDZHba3Og4f+QRE4OA7JmrKEtzF6oyhq0WbmqVsGhqW/BDvzbr1qDFl8UYbOWMzpczBjT
wNlTjLoiZlhkC4PMj46vDSn+r/mlHlJ85SxS+YTTIGOIQpIMNxrl9+AgpwZChF6oTnQGKDqBWra0
kFNhfB/ocmpQu52oQhbDQl8qkzoawxjWb6A4yju8JRMvkE4x56dpSkZ5Tfgzhjtw+0zy7UOFTbGQ
0/TL36PmKVChYflWHzUOSE+oryb5VkNBLGKm4uFmbu1Z4zRnIq81YKUbcy9bzwf21A3iHqZzxMIz
hNsPMGy7uySIqJYVK89Q+2Ra/vrIjdCTN6UEF7E1JNrbnmDmiZg+BWYjJ/ULhS1TmLBlXoS+bVe4
IF35vL2b3ql1foATccbPnRVrHDsJf02XYOOmiRohWFN5WYjjCOEAsuQMKgqzbGC3Wab7IgjiVOrq
z80rqINuXrLAqAqPgZhLq8MzcI5M3Nqpky8MHKs3DE2+QiMqGCe+N5ryeKbAc2p9disiIkSIvOT+
tBVaiswMPGb6W0ULHvUHZPPn9vRzPFd3Tda/x6VXzGEtnB92QfynrYUnqosk44GPXPynuN14iNNV
K5QK6/dKbdEtSF2kcyZl/Q3NfvGXjcNQwjHcJCWJu5/CXNJMvUlbckLN1i2GgYQ43oMZ5RmE6tiv
7h1FLex3kxLEEwF/oCL7PSuvYEJZZsb96Vmpagr7nrbj9WNfpfNQuxElZUJpWke/x9LK+dSNFqGN
Hb1dQfezUV4bF0HBuQqL8BecDYI9CKbTLVUNaMUFZywj6CkbVgtYpndBJWgPRmF2eDD6LwFkwhwS
oUaZl/4cMETKnfJ3korTxAhqIi5EFLhl/DNrByO76Pq9pX7pjNOXH8qdVfrKwtwcWpTS5G4NMcEW
qQykuwG4dV7mlCT7RwAqN7PDFUph2aQA5xs/Olyclj5vG9nH0wG6taPG/OqA9ZhnYKGkMbzmOAxD
aGNgoVojn/2vvN+i8oMplOAM6TGoqBcIglP90UxKYO8jLf2svXrBGt+HVjL6ckwOLtXvHElPuItM
7dk/hk3iwUV99tmXnsyrXSE8ZzKHuEq1JMBWbQftZc0UzxYg8CuvArZUye2qsk3bGYrgf6WQNvuI
/OPr103KEvTRknz0r4S9NPba9vys9FL15gUwXNSF+Cmci7GFyFo6XiIg0d2UOEbziLckwhb6WF6Y
19Atly2ftsaQUvxSqj93BEO+fTZG687aYR2nu8KUEGOJQpOtDU6/OwhOIUVcwR0k/a6E0fR7ezCs
B0J+fW4FuI/h7eD3jmbYRi6RtJap+hLAPKAWuuEwFoNf2WWa/RRCytG7ZhUJ1pEELRgAbVdywZT4
KsqOwHAr0oEoUQRRfCI3uBUxsnTNosQGIelPyORiHGE9geyy/6B9BH/8njLTseds3hHRtyN5gfIc
ajSVHG1KP8gCjEZdu29F8LuiY4RqLz71YO0Aeb7RmxFq4nw3TTRWZ8IAGeEKNZG+h+oSR3YH0qlR
5cCvggwqsQMblTMbYux8gDkepjFJuDqaTyOCL2W+RKiWLRvuJPLC1dnXZjHQ/XlrkshxjWKTWmJf
IEegza0CjVKJbmmAbdUC58Pcjyp8WXP5727xaRLx3VkgKMjntEjcy8MgrrTjpjkgiqQMwlK/4xm2
9SiywaxtWbUb5YmGl5wnBC3O7TzZFU5C/3OuFYjOJscyHAkJleMfLHnZunZQ5vf0K060PMczQyQs
1EE4ZjcpOCBfjpxyjtUOtCrOmx9Rx73t6ZQ5VQf3bZkkDqIKhJ2iN0sssX+5QVZPd6AomaGy1VhT
BVo8pHhcgoflDcyEC+w/no+jW0VOBDV4tpqlHnI+4AYtsO1cMAQLC/9ucb8/4yto8lU/dNqzyd+i
Nv+kBebw0B5kwN8SBAApiC64vaAPBysZDj5PK5jEzxdOmE1czlaQCZ91rNlaZ3jVm1nOJ3trTASI
16rxxGTEOKDJOIq8DlPsk3Cx/mtUUVU/8Tt05gJBiOIOk4pCPxU4Et2rjsvuqY6vkBnIFhw3yauu
THG5UvOQCS6rXzjEsCgAfpFub7KtWLZbWdH4/AVyAs6PET14RliWltpfb6cgGiTzgmq/nscj/ZuL
/WZyeH1rcZcrvf24TVuVdEnJA/aRCKoJprSrb37S9QKNc/vDKuSRj3Zdo9MvutSTO0C70cCg1ftN
PsxGZf0Hdv+BINQVSesSV4/Hv+l2e8iAw3fixLnentvsrsII5EWCf3dUJJ9WTKW3e6S5mblckJ+5
eplPeg5ISCMDBIwh2g/NKfuP/WlPy9evu1h7HByzocf5/QDnyP0sowSIw5ppaS0BtFcm1IvC8arm
J7kdpi9o5S1bvEzwKRmtghBMUnMWl5diqKCwjkdSJ/LZUy1CAwN+cooMztLosoSMUUdpaT0etDyL
+IXpE0tZMOsfUXeehN/4q/8BSiFNoNang/KivRTRSupVV+erLT5h6tpiR8UPelXiJaNnNZuGQSWK
9dP0FxYnPhIwquBy6F4WHWRiUSA+yEqqKBV0p+JJp0TNuWVqi9JSE8hVQ1peLK+OaKL4aitccULM
MHOs0lYb0sNL4t+YD8mhKy08TYAatoymWUSHBTINQcgDLt+GUcuMXZajnUlHzxp8IGPYoQqF1JNn
p2S8uXG/WnFfAZ2PACdO1YvtTbTG/xD6eWLunhD/wdDQDZD0qvNXVH3WfyHYynsvRGtNALcnunxF
brF++ZfSKNvCz+SIU8QdLjny/paJVGBJ4gPxTs2zhXuOZIAjfdEIMFAfWcDrjdrjZdybS3bhU1/k
2d0L2kxJaotLhwWrCji+xBDjVh36ddNT361xVd2yb6MPPCDyCAVRODYUPlY29HSWta+x4EZjUXel
UCvtgBOSuavL3h6nmIOyCDBbeo6oJiOsj0QbSwzy5GVOY2BRt+3XiI+/jTCNqoLI4+ZRtooGafsk
ZlJGn6AgMCUxpmkpmUk2OeXUDXrYKhsPPUJAnwVY98G3QzuEsEZZKp88VAfipwT+B2c4MUWcXZT0
b92WxieZef9nwKwrUHUk2AGZxESRSRzkR0PuUc8644TGmnJvMQfmR+hbE+7p+1hRYF2VeUUz2hmv
bXZI+LjtM/5zBeBu9KED16jBYqEmZLkZkLB6W/89+Ck+4pOxDJKC6Qf8rfGv7eBK+iFnSlKGE1RU
rlS2ykLqsZCl+sYOGsoZRhER457xG+A6XNMBKD3c20wVmBSf2KAoYsArqHJo/DM++yUs14CsCEVN
Mh1pjQtGoOr4i0yngp2/IFqmPJJqBy5os+7ee9OgjWkwJPFhyeswkIZ+g105Fq7uavl+6gk7/KBA
7EGJ+ABXO0WCOzuz/haCwcPVF2lVRKupz0VEE/vUxTbyXClLq3a7CDJxBXRJsirNyvq+RvSmfVW7
ih7cGd88SMCC4YuuTIOY25Ze/+99rkMcmFn6gNLx6GrKiTSsAlO5K9Vm82pqMiZO3pn6cRLlP1OQ
TXHjGycotYQ2zfT7FYZ/w4olYQ0gskgAst7OPJwPy75tQWDBqQpH/y2UQi9Wg6xt4KhP2Kq7vtCa
TkZRrG34OJ8IPS5f73X9yp+4O9FMq57A4bINCJwEkD2yoUHluSoeUsU8AFTJ63wslc3Zwp4IWnZx
GovcmFpmTxbZiie4ysi8njN/EGHii3Ao+zGGWacqfYZ3MJaRck7SdrM8fExpLhGjPF6ykK4xNXKG
1thT8ZrPqJwu5N/0GntUcxHn6Dj2OMK4MOdK8SclCzcfr4ccelIxjOp/+wxw8YjWpzTygbJw4APk
RekDjNK+zV+WKUmT2EWoECP2KMua7hBc7wTDvyZsTjQRvZqBgw8jUgEyvlYq7b37+aaQznAWuBbo
A1xiE7G9bJZ8PmmI8GUzRxC8zs+gsDqkTEJue+EvdJBdlVb7jOv32AUuS4XBDo4bVSlcqgDhn2Xf
HEBVF4IkXaGLcMaoDax9rQ3NhiPiHJ3VF5OXBgkj43PGnXPeraYZ6Q1dVt0mTl/A/KOmJNO5Jz4W
PSWX3l2oPuUUafvxxi+qS3glCsXuXNHZdNWNHLEqZcliO+S9HSfM0sm92fVAfls8Xd97sPC8yCF4
9sMU5UgqrkuhtrEmeAo7JnwCnBTdPUe3sv0PG8c0wewpq6PueTTtSYnTp2m3N/7ZpN/ZLvf9Z6Rm
pThFcJjU1Q5q5kXJ5GqBotTZnUPCTPfvh7l5BpUVOnShxMEONws7kMF3FPyTUANAJovcgS9WJi9v
605JE2GXzgKzsvN6KfnBGpUFbahOgEX5ex/Ymr3+eDv63fVuNdlXanhOLgFuAZScE3znogTarSJa
zWskuFcZ0dmwXl7JEueOSpj7iJS4wXcz+FcB2cDmlPvMfmHnR6D7rSVs2c7RgEB7f6IXfb1CQ4FJ
sx+TgtO1Xm/WyQD6o2nAP0GgJBOy3s+yf6CRs0DX2sWKEHZFHCcR17xA5c7yN1LuPTV/FQnBho2X
kutLdxkbtMzL5IFoAMMns5IfCPnpx4yBWSbIqFIx3AzNV9nQbFtn0z8UgHmpwmArrPfSuTFBtsMW
5aUMcLVOUJtKdfWWm+y4CwEKmqVyasHhiHH1MjRY5s/1dnj4o3YpavTM49WDmom8gSR9jU8iLaX1
WmeOsEf5Y22T4fnwCoL3wtfnwiLCPYuCZcPq2QPm2b/eF2ozXdjdqlLx5DASYN4WwIxHmqAYxd7s
KvNyckluNAM7JJnrYD1Wa5GbFcLIZbaQk8pXIlQquUDYrZcTWtdhO4FHqm0G5/yszh5kmYGqtvdR
E59M2QCALPtVJbVqdcu85ostYhi0XWN2S/Aqdy2NT5i1abSJqM2V2Yt+u6doPnBwcCadQF6G0SLV
V37OLn6GWqJkRxata54kWJqusRwtqqSaKFVZI9QGugbMfRr1QFL9C/vgwOHBeJ3MznhhB1Pm/iy4
Ta+Ah1XG/s0Sh8fsObWt6tuTJmkwBdJNxj/ji0ierGdw3K7Enx/5F1j65xN+vCHsmuIeyc6b7bAv
WifUTq7DtO1sO6q5ZxMRZdm0AHhDnN/tHj7qkfDqOvQseAYytd7m1RkeNailM/Hwjj8TQ84o/fOr
BytCHFQe+75lSxY1Amr3Vys6k4/DuykMZYGG9mcSs607o9qNcMigUMlZ/oonmgO602/pVT4RArzW
UBMVuezXmBa442Vy63ZhwCF5A5/OVbkJnF0Wnu4Eyi2Qm5GB3NYk0bkQKDISjWTZ8j3A4iEG52s1
PL2QKrZuGAn8vR/Mnh9lMgqNYXeM3l6e6cuiDrwOQi+HRpFHFgqV98QI+qM/k56u+50VgkIrlciV
sGF1jSKHp6LDhvl1JwMAMp2IdX8wl84vh9CcA5ztlUirPN4rar55aOCcHMpq4DQ+sxlsJMe26pzq
P6lECOMpgn4lRw5m0h/d1Gvm8qXS8Z9Dz3uHA3yJWoGlw+JOcphdwUymiIYkZnh3tDDLPqM4HYSm
5Lqemk2DJwMeQtDud3FEPd2uL28wELb7wNRGBgdsgbDzdCHe9+vD76vkaCcoPZzkhj8J94M0NEnv
ozgA0HhIwVD67of1+iwPmUdJpd8m4zqNWrtSLwrCkAlEBiKd30TTXuq7zNL/a+qTTDVQwPkqOs+U
ueM6+22l8a3XHlTYwOUXaCyYhbieX/dtIzZZ6K3TuVhtJ9txRrz+O2QDmGSyx47JpYOSwHlCpA4d
0I+JVOEhiD+NllgDEZx4afq/EFiQxfr70QSG/VbNDynZ3r+m+yDXWIJOSKimmdHNtdR9pYveyBMj
HGBGbIMRzWRAaUtn5cK1OwLTKVAbMPZArkUQar53hahdQCsGJ1tDwd6P8Z0XEDLnTK3O6tNTRdil
MteAN3/u8lUGM7fdp5ZlP4cOV4F89uHKRkcrQYXRylsC/xbQkat0lREDp0TlOcuqDDPJElZvOj71
LogeqE85CXJGVRZmyPIVFRzA14zpdHkZw80xmQrVUl9Acs+4T3Oynzv2FOozE4DQkjps/T52D41e
IrI1DRM6UCu7eTtchpBK8TAhQ2Tk0Oh4d/j1Aqete8C6/bR4rcLBXFcd66JKCbAbTwf8BWVT8k6E
rZ/h82IMJ5awo4nf4nLmunMSEs45U+hb0UCY+3qb6HmrspZYRfLxw8LRtW1z4SrXWTwaOMbAtRwU
QWiIeREZ77XUQ/Vzl8N9ub2PguqvX/ckwKiM0whEgKDcpie7nuCfDbGF/YawOnuyr3nvHhzaxmRW
IPxHWwIxXTLpbpQ2E2Pkh3u9CMrk7wwDoix6Si3xWPmueoouyt+nzans0DT/8ckLJx+gT7fwFpT6
JhK5urGOtW6qt2cQfNi6QVIIAziU55SdY9QNIShDrOdQXGhE+LnrN+SHNNBc8/VaHb7zEjtkEiWM
EgizfXSSLC+60uUWeEOORsscBa64T32kXCzkHukkjcJHuWZpeGGdhv5jENmKBr38MGxJlK2IO4Ce
AXRAkZJdNnCZ5XLZ9xxfRLh2o3uasx40YdbD9OfzW6TWEoAO2p/fe3sAltM532TqAQ2CYZAd8OUp
lYGhmnw7DQVimoWXwx2eGGn7+Cn5WSMF+O3n+iRW7KUMfaxRYUk+haAK8jDixN0ZxSlhGMXB9OPm
vRZkCiipjkKheM41bgirak0/LExTRJ5UW2fu9FKo+DmTWWiERfPsD6qob4q9PhEz2aMUxnkaQEUr
JEIBuckDapxNVboo8N2rjmxhsAdnWhtkVtby326V5uZsfgUsr9Egi5iVk+FIn5vr2V1qKVCbr+cd
Vb11LouGQO0NQ0JlwlD/q2CuxDgaGn9YO2s+6YmWck/+8UQDagMF9TCGTDYpWY6pZTVtdKo1a5vf
bRvsIlc43Gn07plLZrskIFamPdIE44Ua1kQb2sEXme/QBh4upq/jGuIACqRkOm5NM9Xl/EDk8Mwn
y2p6i+3MNjOv4XmNIKQkFYjK9L8RBPk/F+jm5eKWvpT+1jmsxl6/TV79B/h2Zm5IwEubP4OaLUWL
K7OxFETigJQA9hg2jcvv7RNwTbR7CCNF6DgMgmxecFS4wxE4MG67Vm7VEWsATSXt9iyJJTKWDvMi
XOZC2opnGtNbgzYTRl38Gj3jG3E0vJB1hkDYNTvbkjJVb560sI62ZyDjL2qgAMBK4hFzGGFpPkUP
4OA9+JR9XrVWu79YRuxrgzLfu65uBwzFBZ9M3VHSOqevBbcLMFlUogaN+l+l4QfPUdhtJj1OcTHF
P1xTc592iNAnvsZEvNbd4mfgJ5nNay83eb1EjNpbL7ixBlVkEMT1Lls2wgLpsJ3u42r370f42Jou
I0JceADBtZaslML5DBoLX9+wvjN4LPK51idRYSocZTQ88U30D4mNkLyOEYv36i7V7SAtye87cmBy
QaxwdAh/0AV9eamzMku5PU3W3l6QhEZiXndFI5sd6NpXyb2iwkcvvBt4dzm1tC1LT9EYeY42cQay
dExz3CBpqDYC9h+Nwzo4cuaj8mgy2hw+jzxJZGvwzJAecNqnIvhydQrR63f/BozMJnjKlEVHfZms
C9N5pW1jH/Whh0gPRUT2Js4/sjwi9Iu/Kcdy1OXznCNAUxYzeJ9Nqa1bDA7aW/aBcqKPTNM70zio
kwnZpuW+bjiOHE4Cb15LRgvFBLeYkgXUJEk0w/DVeTVhBWiKxfHeo16GjfDrZxqZyA9uvgLl/3wG
i05VHtQDR27hLdSLy0l/U1EhHUtOkwbuZ33gBTF/p2WcEG7YWp4L/YOT8b3x+BcYWBlS8qSaWraP
rqx+3Ekqznr7MeeYpYS87N8lg7H3Oie08J2Vfp0h3fm7l3wJ3nlmx7h8pUTzBRrrXK6HehR+xGRR
/NDzfrofqjRU8GBsXQP9XYmNiG2l+Vc2vOPfM5Cwrfz6K4qfWGfDz9Nq9MYA/QGl/aiRs42tT4DC
WJMD8T6CL4qqSkwBB+ZYwxfRHOz3OkYe3IbbH4FT3RfFtnXwqJ8n4mkr8cz3Ki8aY1RbNlkTsfT+
hM7ikfRbUimkYXjwc41VhkrlJUMvCCnJwwnft+1cccgEmA+hbkZeXc99akBgxNegUgjZYeTeWRfi
MqCByKg4YyPdQjGZ6/By+CnAXVoE+Sr1dBjegN9jts3pCHJnKEcai5lsd10H7outcVUqc5av+R+R
ExohDSpm07e5JTSpg1a/TR+PiSSZtOn66IOwiNqdj9df4fgxUn/SfrPRTuC5Kdr2pcRrO02AV9u0
Xp1qcP+m4uVBR0LUQZX+Ml85ETdaxqmZ9G16PeIoxHtlsSdSSCO5q1UljCZSkXWdCx9alpZtZUa/
6OkIFmLZTPTllMkNDyIXhqJ9+MI0cpHfV9NZI2RBsskI4/++bU6WgujC6fPaz5H8CqSeX5ALfSyp
ejFoZdAGapNFeX1x1O/I8qUIsekP7x100rVdLk0BaAIC0f+3o2H5rpFbJ0y0RYhvyL6W7zIvNRUE
8El1BBJjIsZ/F8FJzFJYRy2aVdb+pk2Gr/cnBc1MM0oPUwZWaO274hs0+5/tDMcD8p7F13nDHoOr
FA3Et1hfGGZH3GPy6FqwUjuqty0+AKbUsv5gOx7/t81WWNAVvw0kg6Z1BfIp2fqwBBPOzDNuuKBk
b7wNY8X7NETjoMN0oZqBwSZbm7ESFxayxtTw31ekV8+ZJC7DWjxNmOcjMRKmimZW7yp4U6aeciP4
NgaIQXxIP+hCvlshDxbddagBEfL7fqBjIhbMmgk9j2Avsu3BisICSlaeVIRjtxkTAM7T12D9fIhP
0+j9dqo3bRrgLCQtmj8neN/sUfkFwSNnLHusXThnEKUkJ1KP5sInbc3b34Gn9mRpHUN+dqFnXV6q
6ol1gD7x/0/q2LrsI2YUZaxjtuZ+feOk3xVAKLbuh1xN+hBJSgLaKy2EeffNnjhVZ9R1i/uOfwuv
AnLochvIVFkEDusxkLmI+Hz7WIkNDcEWChRZYey2yf53tm28JHN08BemCR8+VlV5SbFIxircVHnF
G2ITiirEQlvqOT9yQcsTRsU4KC7M5s1WZba8xF0UbARAVFemOxuCsROjSWBc9AJ5ehh6+zTRwuQE
c+1DhLglCLydI+G/lUwW6KPCg4EvgARt+cDpi8B2W7mSWWp1WB46vo4hMzv+wcqFA/lMn6k6MjPz
1BkXNhmHkGFuzvF3l/QJiaDnIS0FpCESUjK6/8uNR4ddiXzF5XZH7hT0rVTLQ9Bsz6o6CXcorCJ1
n1lZHuHZsJ82foNhFKisQdZ484sM1tq6A25BxB6IuJ32C491OP6odIdCOveTnQC3KFliuwXRsVLT
OhSeJWM+/vznu5MiSb+qZGUgfs9uyodNznqWTu6Mz/k6GnaDi+NqqpuRUrJq0nGi+jU4tYb5CeC5
8AtVTnVdU9v3xEuTsudEAGaNTRu8IocW34gu8IDm1RpSaefiD1RcNuWRF6vJai+sPw66EbeSnj3S
2bKL+Qkh7p0Xd5GqBULK9XhXCn5mJItkT6G8xYq3knovgNWssixTHT93qvpabH1WxciM8OIUgE6H
AwH4sWP9ba7HpD2W97reCepEyf+rT/heufTrrZnYchGVBhn0rtN7c9FuLq5LbfYkLLuztOwJo3h2
Lps/WuZHE+WU9AlMWe/NLXZJAjCkdFM04naIl+28IEF0ff0HoEd3V6XgT1Y7x0AIDcv+pAQLXLOY
GpqfIjFMwCmK4LPO4Cr6bv+uAhe5RARS5F/IM/KFhqezOt7T50lg5Rnm6Df5f3vMW9yLIFZf1o2X
AN1+K0H3jAiq0XEztAFQGXniSZSp0qH8O8oMIGWhNUbbVh370it6KzAi2Mcr228rJGmSHg0qhOG4
jOeDMKFActNzw1YNWJ0dEmNBfXbhWGanoXMju8CutFUeMdCwn19WkNTzgztWOoD8WeXofpH5BNg/
1gPzuUWtnTeVMXUwZWdteSetL6N0qsKM2QjxoZBPL7Hj8Ru+3N/RcuS7d+dsvMK9xRTJcMPhkyo5
T3hip8urTAx4uiPC+l6d1PJ5NpNJjWRC/gvP52/1Tp6oBt1gemcEj81K7OpiJMRlEanekLLCi0N1
fbqiEbfQyN9+wNT77SfAKxMdLxOZFDRwyJppzaDvgVRqZOLd/Mum1grnzGRoNnkFDIbyQ+u6iMga
hHwI6HQAfFPebLFBySauQVvXt3GdpV14schRJ4U2XAnQIJ1r6aLZ5YlERWUaLnbY840tnWZPHMqJ
ehhpKNuPV5TEN+ziuecGx1VcACiBATgj+M8/HKkdyOUK5fX+CzkSoTgq/kuhsCzvAv2+bAdeVz8R
eYgUh2fpULazeO76/fpTZrz+kaYYd71PjFcVGeJBmtQNWEtmFUuqPQuBNWw3WbYTj+hAePNHOvYd
gTH2+RxdxK0QfVKzP2vsBIYNi6WxdWR34koJh0Z+8tb//mOtRNiXljjAbAA4ybqJ5z30+S/XVbtF
mRhFosxRj1O7VD1y14bB2ymEz3pWqcGoVfN1iJYOANx3oV8u+PfAEE7Uxs7VxpF2OaHpsSLTyP8b
Na8PSEn872e4fbIv+LPhMJJvFD8OR1XNzbnBZT2lb8OdR+tlyu8w8jLPa2UuTzMNsnWbOqPcqJ0d
HrxkryUF6gAYNKSzuyqs/M4oyczRq9/fbnm+UuaZ35vbdLyKkt6IqcEI7BU3HZp0lkeF+7DTCI2F
MOOfLySTTOnzYz4JsJ/8pQ5HmAc7s3llzLdfKBY6EWyWiQPThjWcdSJaU3cNcvTomf/kT95YN1Vg
78/9jK5XkRkl8diF7nKsbKqE5jbQVKDBTNgtoKOHbos/+M0aziU/PTFEuxUD6v7/Z+xxkpPMTCSf
GJcYd9mPXnGQ1n6+fWhBHXOUc2HrSTW9LmYzvjNZrQLJUxmktLMj0MkW8ZlDqelSyVK/EnS78Srl
S3XNaMPtWRyS8He4OC8nB5AttxjgAWafPd7EqkRR6KhIXawgtEUwG27GCdZDh49vJwqf++l781hB
v9f3PRe5Fv/Z0bPq2BFMjVGOmjkKUy+KWuOFHUcq79cFuf8Z3+MUgvRoqM1zmT+e6cYAI3fw1bYP
Z2P78v/G5cZukpdsiJ6sdzU7gmIE82+jqQMfoOaHOEv5S2v09v08Qx+V1R3Y8ACnHGz0JFRGf9xS
ijDwTFQ9QG4ixr0vVodijodLxjjP
`pragma protect end_protected
